magic
tech sky130A
magscale 1 2
timestamp 1647557548
<< viali >>
rect 29009 49317 29043 49351
rect 6561 49249 6595 49283
rect 7113 49249 7147 49283
rect 9413 49249 9447 49283
rect 12725 49249 12759 49283
rect 16681 49249 16715 49283
rect 16957 49249 16991 49283
rect 22569 49249 22603 49283
rect 29745 49249 29779 49283
rect 30941 49249 30975 49283
rect 43177 49249 43211 49283
rect 45569 49249 45603 49283
rect 1869 49181 1903 49215
rect 4261 49181 4295 49215
rect 5089 49181 5123 49215
rect 8953 49181 8987 49215
rect 11989 49181 12023 49215
rect 13001 49181 13035 49215
rect 14565 49181 14599 49215
rect 15393 49181 15427 49215
rect 18153 49181 18187 49215
rect 19441 49181 19475 49215
rect 20085 49181 20119 49215
rect 21281 49181 21315 49215
rect 21833 49181 21867 49215
rect 24593 49181 24627 49215
rect 25973 49181 26007 49215
rect 27445 49181 27479 49215
rect 28273 49181 28307 49215
rect 28825 49181 28859 49215
rect 33057 49181 33091 49215
rect 33793 49181 33827 49215
rect 35541 49181 35575 49215
rect 36185 49181 36219 49215
rect 38209 49181 38243 49215
rect 40233 49181 40267 49215
rect 42625 49181 42659 49215
rect 45017 49181 45051 49215
rect 47777 49181 47811 49215
rect 2789 49113 2823 49147
rect 2973 49113 3007 49147
rect 6745 49113 6779 49147
rect 9137 49113 9171 49147
rect 19625 49113 19659 49147
rect 22017 49113 22051 49147
rect 27629 49113 27663 49147
rect 29929 49113 29963 49147
rect 40785 49113 40819 49147
rect 41521 49113 41555 49147
rect 42809 49113 42843 49147
rect 45201 49113 45235 49147
rect 1961 49045 1995 49079
rect 4537 49045 4571 49079
rect 5273 49045 5307 49079
rect 12081 49045 12115 49079
rect 14657 49045 14691 49079
rect 15209 49045 15243 49079
rect 20269 49045 20303 49079
rect 21097 49045 21131 49079
rect 24409 49045 24443 49079
rect 26065 49045 26099 49079
rect 32229 49045 32263 49079
rect 38301 49045 38335 49079
rect 40877 49045 40911 49079
rect 41613 49045 41647 49079
rect 47869 49045 47903 49079
rect 41797 48841 41831 48875
rect 3525 48773 3559 48807
rect 9321 48773 9355 48807
rect 35081 48773 35115 48807
rect 36737 48773 36771 48807
rect 44741 48773 44775 48807
rect 47777 48773 47811 48807
rect 19165 48705 19199 48739
rect 21281 48705 21315 48739
rect 32137 48705 32171 48739
rect 34897 48705 34931 48739
rect 41705 48705 41739 48739
rect 1685 48637 1719 48671
rect 1869 48637 1903 48671
rect 3985 48637 4019 48671
rect 4169 48637 4203 48671
rect 5641 48637 5675 48671
rect 6377 48637 6411 48671
rect 6561 48637 6595 48671
rect 7757 48637 7791 48671
rect 9137 48637 9171 48671
rect 9689 48637 9723 48671
rect 12449 48637 12483 48671
rect 12633 48637 12667 48671
rect 12909 48637 12943 48671
rect 16129 48637 16163 48671
rect 16681 48637 16715 48671
rect 16865 48637 16899 48671
rect 17141 48637 17175 48671
rect 22017 48637 22051 48671
rect 22477 48637 22511 48671
rect 22661 48637 22695 48671
rect 23489 48637 23523 48671
rect 26433 48637 26467 48671
rect 27077 48637 27111 48671
rect 27261 48637 27295 48671
rect 27813 48637 27847 48671
rect 29377 48637 29411 48671
rect 29561 48637 29595 48671
rect 29837 48637 29871 48671
rect 32321 48637 32355 48671
rect 33149 48637 33183 48671
rect 38761 48637 38795 48671
rect 39221 48637 39255 48671
rect 39405 48637 39439 48671
rect 40049 48637 40083 48671
rect 42901 48637 42935 48671
rect 43085 48637 43119 48671
rect 45201 48637 45235 48671
rect 45385 48637 45419 48671
rect 45753 48637 45787 48671
rect 11713 48501 11747 48535
rect 14933 48501 14967 48535
rect 18981 48501 19015 48535
rect 20453 48501 20487 48535
rect 24961 48501 24995 48535
rect 25789 48501 25823 48535
rect 47869 48501 47903 48535
rect 12725 48297 12759 48331
rect 13461 48297 13495 48331
rect 22937 48297 22971 48331
rect 29653 48297 29687 48331
rect 34805 48297 34839 48331
rect 39957 48297 39991 48331
rect 7389 48229 7423 48263
rect 8033 48229 8067 48263
rect 30665 48229 30699 48263
rect 44097 48229 44131 48263
rect 1869 48161 1903 48195
rect 4537 48161 4571 48195
rect 5641 48161 5675 48195
rect 9229 48161 9263 48195
rect 9873 48161 9907 48195
rect 14473 48161 14507 48195
rect 15209 48161 15243 48195
rect 16865 48161 16899 48195
rect 18061 48161 18095 48195
rect 20269 48161 20303 48195
rect 20729 48161 20763 48195
rect 24409 48161 24443 48195
rect 25053 48161 25087 48195
rect 26709 48161 26743 48195
rect 27169 48161 27203 48195
rect 31309 48161 31343 48195
rect 32229 48161 32263 48195
rect 35449 48161 35483 48195
rect 36277 48161 36311 48195
rect 42533 48161 42567 48195
rect 46305 48161 46339 48195
rect 46857 48161 46891 48195
rect 1409 48093 1443 48127
rect 3801 48093 3835 48127
rect 7297 48093 7331 48127
rect 7941 48093 7975 48127
rect 13369 48093 13403 48127
rect 22845 48093 22879 48127
rect 23673 48093 23707 48127
rect 29561 48093 29595 48127
rect 30573 48093 30607 48127
rect 33609 48093 33643 48127
rect 34713 48093 34747 48127
rect 39865 48093 39899 48127
rect 40969 48093 41003 48127
rect 41429 48093 41463 48127
rect 43913 48093 43947 48127
rect 45017 48093 45051 48127
rect 1593 48025 1627 48059
rect 4721 48025 4755 48059
rect 10057 48025 10091 48059
rect 11713 48025 11747 48059
rect 14657 48025 14691 48059
rect 17049 48025 17083 48059
rect 20453 48025 20487 48059
rect 23765 48025 23799 48059
rect 24593 48025 24627 48059
rect 26893 48025 26927 48059
rect 31493 48025 31527 48059
rect 35633 48025 35667 48059
rect 41613 48025 41647 48059
rect 46489 48025 46523 48059
rect 3985 47957 4019 47991
rect 33701 47957 33735 47991
rect 45201 47957 45235 47991
rect 4353 47753 4387 47787
rect 4997 47753 5031 47787
rect 9873 47753 9907 47787
rect 10517 47753 10551 47787
rect 14381 47753 14415 47787
rect 16773 47753 16807 47787
rect 17417 47753 17451 47787
rect 20269 47753 20303 47787
rect 22293 47753 22327 47787
rect 26341 47753 26375 47787
rect 27445 47753 27479 47787
rect 31125 47753 31159 47787
rect 32505 47753 32539 47787
rect 41797 47753 41831 47787
rect 5641 47685 5675 47719
rect 33701 47685 33735 47719
rect 35909 47685 35943 47719
rect 43913 47685 43947 47719
rect 47777 47685 47811 47719
rect 4261 47617 4295 47651
rect 4905 47617 4939 47651
rect 8861 47617 8895 47651
rect 9781 47617 9815 47651
rect 10425 47617 10459 47651
rect 14289 47617 14323 47651
rect 16681 47617 16715 47651
rect 17325 47617 17359 47651
rect 20177 47617 20211 47651
rect 20821 47617 20855 47651
rect 22201 47617 22235 47651
rect 26249 47617 26283 47651
rect 27353 47617 27387 47651
rect 27997 47617 28031 47651
rect 30481 47617 30515 47651
rect 31033 47617 31067 47651
rect 32413 47617 32447 47651
rect 33517 47617 33551 47651
rect 35817 47617 35851 47651
rect 41245 47617 41279 47651
rect 41705 47617 41739 47651
rect 42533 47617 42567 47651
rect 43637 47617 43671 47651
rect 1961 47549 1995 47583
rect 2145 47549 2179 47583
rect 3157 47549 3191 47583
rect 6377 47549 6411 47583
rect 6561 47549 6595 47583
rect 6929 47549 6963 47583
rect 28181 47549 28215 47583
rect 28457 47549 28491 47583
rect 34713 47549 34747 47583
rect 43085 47549 43119 47583
rect 45109 47549 45143 47583
rect 45293 47549 45327 47583
rect 46581 47549 46615 47583
rect 5733 47413 5767 47447
rect 20913 47413 20947 47447
rect 47869 47413 47903 47447
rect 3893 47209 3927 47243
rect 4813 47209 4847 47243
rect 5549 47209 5583 47243
rect 6285 47209 6319 47243
rect 7021 47209 7055 47243
rect 7849 47209 7883 47243
rect 27905 47209 27939 47243
rect 45109 47209 45143 47243
rect 1409 47073 1443 47107
rect 1869 47073 1903 47107
rect 20545 47073 20579 47107
rect 43637 47073 43671 47107
rect 46305 47073 46339 47107
rect 46765 47073 46799 47107
rect 3801 47005 3835 47039
rect 4721 47005 4755 47039
rect 6193 47005 6227 47039
rect 7757 47005 7791 47039
rect 20361 47005 20395 47039
rect 27813 47005 27847 47039
rect 41613 47005 41647 47039
rect 43269 47005 43303 47039
rect 45017 47005 45051 47039
rect 45661 47005 45695 47039
rect 1593 46937 1627 46971
rect 22201 46937 22235 46971
rect 42349 46937 42383 46971
rect 46489 46937 46523 46971
rect 45753 46869 45787 46903
rect 2881 46665 2915 46699
rect 44097 46665 44131 46699
rect 45385 46597 45419 46631
rect 47041 46597 47075 46631
rect 47961 46597 47995 46631
rect 1593 46529 1627 46563
rect 2053 46529 2087 46563
rect 2789 46529 2823 46563
rect 3617 46529 3651 46563
rect 4261 46529 4295 46563
rect 5365 46529 5399 46563
rect 42625 46529 42659 46563
rect 44005 46529 44039 46563
rect 42809 46461 42843 46495
rect 45201 46461 45235 46495
rect 2237 46325 2271 46359
rect 48053 46325 48087 46359
rect 2421 46121 2455 46155
rect 3985 46121 4019 46155
rect 42441 46121 42475 46155
rect 43821 46121 43855 46155
rect 44465 46121 44499 46155
rect 45109 46121 45143 46155
rect 45753 46121 45787 46155
rect 48145 45985 48179 46019
rect 1409 45917 1443 45951
rect 2329 45917 2363 45951
rect 3157 45917 3191 45951
rect 42257 45917 42291 45951
rect 45017 45917 45051 45951
rect 45661 45917 45695 45951
rect 46305 45917 46339 45951
rect 46489 45849 46523 45883
rect 1593 45781 1627 45815
rect 41981 45781 42015 45815
rect 47685 45509 47719 45543
rect 1777 45441 1811 45475
rect 44097 45441 44131 45475
rect 44741 45441 44775 45475
rect 47593 45441 47627 45475
rect 1961 45373 1995 45407
rect 2789 45373 2823 45407
rect 45201 45373 45235 45407
rect 45385 45373 45419 45407
rect 46857 45373 46891 45407
rect 45201 45033 45235 45067
rect 45753 45033 45787 45067
rect 2789 44897 2823 44931
rect 46305 44897 46339 44931
rect 48145 44897 48179 44931
rect 1409 44829 1443 44863
rect 45661 44829 45695 44863
rect 1593 44761 1627 44795
rect 46489 44761 46523 44795
rect 2789 44489 2823 44523
rect 3433 44489 3467 44523
rect 46949 44489 46983 44523
rect 47685 44489 47719 44523
rect 1869 44353 1903 44387
rect 2697 44353 2731 44387
rect 3341 44353 3375 44387
rect 45293 44353 45327 44387
rect 46397 44353 46431 44387
rect 46857 44353 46891 44387
rect 47593 44353 47627 44387
rect 2145 44149 2179 44183
rect 2881 43945 2915 43979
rect 46765 43945 46799 43979
rect 47409 43877 47443 43911
rect 27721 43809 27755 43843
rect 27261 43741 27295 43775
rect 47869 43741 47903 43775
rect 1869 43673 1903 43707
rect 1961 43605 1995 43639
rect 48053 43605 48087 43639
rect 47961 43265 47995 43299
rect 47041 43061 47075 43095
rect 48053 43061 48087 43095
rect 46305 42721 46339 42755
rect 48145 42721 48179 42755
rect 46489 42585 46523 42619
rect 47593 42245 47627 42279
rect 22753 42177 22787 42211
rect 22937 42177 22971 42211
rect 23029 42177 23063 42211
rect 47869 42177 47903 42211
rect 2053 41973 2087 42007
rect 22569 41973 22603 42007
rect 1409 41633 1443 41667
rect 1869 41633 1903 41667
rect 46305 41633 46339 41667
rect 19257 41565 19291 41599
rect 21281 41565 21315 41599
rect 23397 41565 23431 41599
rect 23489 41565 23523 41599
rect 23581 41565 23615 41599
rect 23765 41565 23799 41599
rect 1593 41497 1627 41531
rect 19524 41497 19558 41531
rect 21548 41497 21582 41531
rect 46489 41497 46523 41531
rect 48145 41497 48179 41531
rect 20637 41429 20671 41463
rect 22661 41429 22695 41463
rect 23121 41429 23155 41463
rect 2605 41225 2639 41259
rect 18889 41225 18923 41259
rect 21833 41225 21867 41259
rect 46765 41225 46799 41259
rect 23480 41157 23514 41191
rect 1869 41089 1903 41123
rect 2513 41089 2547 41123
rect 19165 41089 19199 41123
rect 19257 41089 19291 41123
rect 19349 41089 19383 41123
rect 19533 41089 19567 41123
rect 20177 41089 20211 41123
rect 20361 41089 20395 41123
rect 20453 41089 20487 41123
rect 22109 41089 22143 41123
rect 22201 41089 22235 41123
rect 22293 41089 22327 41123
rect 22477 41089 22511 41123
rect 46673 41089 46707 41123
rect 47777 41089 47811 41123
rect 19993 41021 20027 41055
rect 23213 41021 23247 41055
rect 2053 40953 2087 40987
rect 24593 40885 24627 40919
rect 21649 40681 21683 40715
rect 24501 40545 24535 40579
rect 47317 40545 47351 40579
rect 1409 40477 1443 40511
rect 19625 40477 19659 40511
rect 19901 40477 19935 40511
rect 21833 40477 21867 40511
rect 22109 40477 22143 40511
rect 22753 40477 22787 40511
rect 22937 40477 22971 40511
rect 23029 40477 23063 40511
rect 47593 40477 47627 40511
rect 22569 40409 22603 40443
rect 24746 40409 24780 40443
rect 1593 40341 1627 40375
rect 19441 40341 19475 40375
rect 19809 40341 19843 40375
rect 22017 40341 22051 40375
rect 25881 40341 25915 40375
rect 20453 40137 20487 40171
rect 24593 40137 24627 40171
rect 26065 40137 26099 40171
rect 26985 40137 27019 40171
rect 27353 40069 27387 40103
rect 28181 40069 28215 40103
rect 28365 40069 28399 40103
rect 18429 40001 18463 40035
rect 19329 40001 19363 40035
rect 23009 40001 23043 40035
rect 24869 40001 24903 40035
rect 24961 40001 24995 40035
rect 25053 40001 25087 40035
rect 25237 40001 25271 40035
rect 25881 40001 25915 40035
rect 26157 40001 26191 40035
rect 47593 40001 47627 40035
rect 19073 39933 19107 39967
rect 22753 39933 22787 39967
rect 27445 39933 27479 39967
rect 27537 39933 27571 39967
rect 18613 39865 18647 39899
rect 24133 39797 24167 39831
rect 25697 39797 25731 39831
rect 28549 39797 28583 39831
rect 47041 39797 47075 39831
rect 47685 39797 47719 39831
rect 19257 39593 19291 39627
rect 22661 39593 22695 39627
rect 20821 39457 20855 39491
rect 25053 39457 25087 39491
rect 46305 39457 46339 39491
rect 46489 39457 46523 39491
rect 48145 39457 48179 39491
rect 17325 39389 17359 39423
rect 19533 39389 19567 39423
rect 19625 39389 19659 39423
rect 19717 39389 19751 39423
rect 19901 39389 19935 39423
rect 20545 39389 20579 39423
rect 22937 39389 22971 39423
rect 23029 39389 23063 39423
rect 23121 39389 23155 39423
rect 23305 39389 23339 39423
rect 24777 39389 24811 39423
rect 26249 39389 26283 39423
rect 28641 39389 28675 39423
rect 28733 39389 28767 39423
rect 28825 39389 28859 39423
rect 29009 39389 29043 39423
rect 29561 39389 29595 39423
rect 17570 39321 17604 39355
rect 24869 39321 24903 39355
rect 26494 39321 26528 39355
rect 18705 39253 18739 39287
rect 24409 39253 24443 39287
rect 27629 39253 27663 39287
rect 28365 39253 28399 39287
rect 29745 39253 29779 39287
rect 17417 39049 17451 39083
rect 19809 39049 19843 39083
rect 22937 39049 22971 39083
rect 24409 39049 24443 39083
rect 25697 39049 25731 39083
rect 27813 39049 27847 39083
rect 29929 39049 29963 39083
rect 48053 39049 48087 39083
rect 19441 38981 19475 39015
rect 22845 38981 22879 39015
rect 24041 38981 24075 39015
rect 28794 38981 28828 39015
rect 17693 38913 17727 38947
rect 17785 38913 17819 38947
rect 17877 38913 17911 38947
rect 18061 38913 18095 38947
rect 18521 38913 18555 38947
rect 19625 38913 19659 38947
rect 19901 38913 19935 38947
rect 24225 38913 24259 38947
rect 24869 38913 24903 38947
rect 25973 38913 26007 38947
rect 26065 38913 26099 38947
rect 26157 38913 26191 38947
rect 26341 38913 26375 38947
rect 27721 38913 27755 38947
rect 28549 38913 28583 38947
rect 47961 38913 47995 38947
rect 2053 38845 2087 38879
rect 2237 38845 2271 38879
rect 2881 38845 2915 38879
rect 24961 38845 24995 38879
rect 27905 38845 27939 38879
rect 18705 38709 18739 38743
rect 24961 38709 24995 38743
rect 25237 38709 25271 38743
rect 27353 38709 27387 38743
rect 47041 38709 47075 38743
rect 2329 38505 2363 38539
rect 23121 38505 23155 38539
rect 23581 38505 23615 38539
rect 24961 38505 24995 38539
rect 30941 38505 30975 38539
rect 17785 38437 17819 38471
rect 19901 38437 19935 38471
rect 23213 38369 23247 38403
rect 29561 38369 29595 38403
rect 46305 38369 46339 38403
rect 48145 38369 48179 38403
rect 17601 38301 17635 38335
rect 22247 38301 22281 38335
rect 22385 38301 22419 38335
rect 22477 38301 22511 38335
rect 22661 38301 22695 38335
rect 23397 38301 23431 38335
rect 24961 38301 24995 38335
rect 25145 38301 25179 38335
rect 27537 38301 27571 38335
rect 27721 38301 27755 38335
rect 28641 38301 28675 38335
rect 28733 38301 28767 38335
rect 28825 38301 28859 38335
rect 29009 38301 29043 38335
rect 18337 38233 18371 38267
rect 19717 38233 19751 38267
rect 23121 38233 23155 38267
rect 28365 38233 28399 38267
rect 29806 38233 29840 38267
rect 46489 38233 46523 38267
rect 18429 38165 18463 38199
rect 22017 38165 22051 38199
rect 25329 38165 25363 38199
rect 27905 38165 27939 38199
rect 3065 37961 3099 37995
rect 23857 37961 23891 37995
rect 24685 37961 24719 37995
rect 25973 37961 26007 37995
rect 46949 37961 46983 37995
rect 22722 37893 22756 37927
rect 24777 37893 24811 37927
rect 1869 37825 1903 37859
rect 2973 37825 3007 37859
rect 18245 37825 18279 37859
rect 18429 37825 18463 37859
rect 20867 37825 20901 37859
rect 20986 37828 21020 37862
rect 21102 37825 21136 37859
rect 21281 37825 21315 37859
rect 25513 37825 25547 37859
rect 25789 37825 25823 37859
rect 29193 37825 29227 37859
rect 29285 37825 29319 37859
rect 29377 37825 29411 37859
rect 29561 37825 29595 37859
rect 46857 37825 46891 37859
rect 47869 37825 47903 37859
rect 22477 37757 22511 37791
rect 24961 37757 24995 37791
rect 25697 37757 25731 37791
rect 1961 37621 1995 37655
rect 18613 37621 18647 37655
rect 20637 37621 20671 37655
rect 24317 37621 24351 37655
rect 25789 37621 25823 37655
rect 28917 37621 28951 37655
rect 48053 37621 48087 37655
rect 19257 37417 19291 37451
rect 23857 37417 23891 37451
rect 27905 37349 27939 37383
rect 1409 37281 1443 37315
rect 19901 37281 19935 37315
rect 24869 37281 24903 37315
rect 25053 37281 25087 37315
rect 29561 37281 29595 37315
rect 1685 37213 1719 37247
rect 7297 37213 7331 37247
rect 17325 37213 17359 37247
rect 19717 37213 19751 37247
rect 21005 37213 21039 37247
rect 21261 37213 21295 37247
rect 23489 37213 23523 37247
rect 24777 37213 24811 37247
rect 29817 37213 29851 37247
rect 46305 37213 46339 37247
rect 17592 37145 17626 37179
rect 19625 37145 19659 37179
rect 23673 37145 23707 37179
rect 27721 37145 27755 37179
rect 46489 37145 46523 37179
rect 48145 37145 48179 37179
rect 7389 37077 7423 37111
rect 18705 37077 18739 37111
rect 22385 37077 22419 37111
rect 24409 37077 24443 37111
rect 30941 37077 30975 37111
rect 24225 36873 24259 36907
rect 25789 36873 25823 36907
rect 29653 36873 29687 36907
rect 47685 36873 47719 36907
rect 7389 36805 7423 36839
rect 20545 36805 20579 36839
rect 23857 36805 23891 36839
rect 18061 36737 18095 36771
rect 18153 36737 18187 36771
rect 18245 36737 18279 36771
rect 18429 36737 18463 36771
rect 19625 36737 19659 36771
rect 19717 36737 19751 36771
rect 24041 36737 24075 36771
rect 25697 36737 25731 36771
rect 27077 36737 27111 36771
rect 27813 36737 27847 36771
rect 28069 36737 28103 36771
rect 29837 36737 29871 36771
rect 30021 36737 30055 36771
rect 30113 36737 30147 36771
rect 47041 36737 47075 36771
rect 47593 36737 47627 36771
rect 7205 36669 7239 36703
rect 8309 36669 8343 36703
rect 19901 36669 19935 36703
rect 25973 36669 26007 36703
rect 20729 36601 20763 36635
rect 2329 36533 2363 36567
rect 17785 36533 17819 36567
rect 19257 36533 19291 36567
rect 25329 36533 25363 36567
rect 27169 36533 27203 36567
rect 29193 36533 29227 36567
rect 8217 36329 8251 36363
rect 17141 36329 17175 36363
rect 17693 36329 17727 36363
rect 19625 36329 19659 36363
rect 24869 36329 24903 36363
rect 26893 36329 26927 36363
rect 21649 36261 21683 36295
rect 22293 36193 22327 36227
rect 2973 36125 3007 36159
rect 6837 36125 6871 36159
rect 17049 36125 17083 36159
rect 17923 36125 17957 36159
rect 18058 36122 18092 36156
rect 18153 36125 18187 36159
rect 18337 36125 18371 36159
rect 19257 36125 19291 36159
rect 19441 36125 19475 36159
rect 20177 36125 20211 36159
rect 20821 36125 20855 36159
rect 22109 36125 22143 36159
rect 24777 36125 24811 36159
rect 27149 36125 27183 36159
rect 27242 36125 27276 36159
rect 27353 36122 27387 36156
rect 27537 36125 27571 36159
rect 47869 36125 47903 36159
rect 7104 36057 7138 36091
rect 21005 36057 21039 36091
rect 23581 36057 23615 36091
rect 25973 36057 26007 36091
rect 26157 36057 26191 36091
rect 3065 35989 3099 36023
rect 20269 35989 20303 36023
rect 21189 35989 21223 36023
rect 22017 35989 22051 36023
rect 23673 35989 23707 36023
rect 26341 35989 26375 36023
rect 48053 35989 48087 36023
rect 7665 35785 7699 35819
rect 25605 35785 25639 35819
rect 25973 35785 26007 35819
rect 28733 35785 28767 35819
rect 2237 35717 2271 35751
rect 17417 35717 17451 35751
rect 20637 35717 20671 35751
rect 24133 35717 24167 35751
rect 24777 35717 24811 35751
rect 26065 35717 26099 35751
rect 2053 35649 2087 35683
rect 7849 35649 7883 35683
rect 17233 35649 17267 35683
rect 18144 35649 18178 35683
rect 20867 35649 20901 35683
rect 20986 35649 21020 35683
rect 21097 35649 21131 35683
rect 21281 35649 21315 35683
rect 21833 35649 21867 35683
rect 22089 35649 22123 35683
rect 23949 35649 23983 35683
rect 24961 35649 24995 35683
rect 27353 35649 27387 35683
rect 27609 35649 27643 35683
rect 2789 35581 2823 35615
rect 17877 35581 17911 35615
rect 26249 35581 26283 35615
rect 19257 35445 19291 35479
rect 23213 35445 23247 35479
rect 25145 35445 25179 35479
rect 47777 35445 47811 35479
rect 15577 35241 15611 35275
rect 24593 35241 24627 35275
rect 26801 35241 26835 35275
rect 28089 35241 28123 35275
rect 20821 35173 20855 35207
rect 22569 35173 22603 35207
rect 1685 35105 1719 35139
rect 11437 35105 11471 35139
rect 13277 35105 13311 35139
rect 19901 35105 19935 35139
rect 23213 35105 23247 35139
rect 24501 35105 24535 35139
rect 25513 35105 25547 35139
rect 25697 35105 25731 35139
rect 32781 35105 32815 35139
rect 46305 35105 46339 35139
rect 48145 35105 48179 35139
rect 1409 35037 1443 35071
rect 15485 35037 15519 35071
rect 17923 35037 17957 35071
rect 18058 35037 18092 35071
rect 18158 35037 18192 35071
rect 18337 35037 18371 35071
rect 19625 35037 19659 35071
rect 20453 35037 20487 35071
rect 21537 35037 21571 35071
rect 21649 35037 21683 35071
rect 21741 35037 21775 35071
rect 21925 35037 21959 35071
rect 24685 35037 24719 35071
rect 25605 35037 25639 35071
rect 27077 35037 27111 35071
rect 27166 35037 27200 35071
rect 27261 35037 27295 35071
rect 27445 35037 27479 35071
rect 32321 35037 32355 35071
rect 11621 34969 11655 35003
rect 19717 34969 19751 35003
rect 20637 34969 20671 35003
rect 22937 34969 22971 35003
rect 24409 34969 24443 35003
rect 25329 34969 25363 35003
rect 27997 34969 28031 35003
rect 32505 34969 32539 35003
rect 46489 34969 46523 35003
rect 17693 34901 17727 34935
rect 19257 34901 19291 34935
rect 21281 34901 21315 34935
rect 23029 34901 23063 34935
rect 24869 34901 24903 34935
rect 25421 34901 25455 34935
rect 11621 34697 11655 34731
rect 19165 34697 19199 34731
rect 19625 34697 19659 34731
rect 23213 34697 23247 34731
rect 25421 34697 25455 34731
rect 26341 34697 26375 34731
rect 33517 34697 33551 34731
rect 18030 34629 18064 34663
rect 21097 34629 21131 34663
rect 31217 34629 31251 34663
rect 36185 34629 36219 34663
rect 11529 34561 11563 34595
rect 17785 34561 17819 34595
rect 19809 34561 19843 34595
rect 21833 34561 21867 34595
rect 22089 34561 22123 34595
rect 25329 34561 25363 34595
rect 26249 34561 26283 34595
rect 26985 34561 27019 34595
rect 27813 34561 27847 34595
rect 28641 34561 28675 34595
rect 29331 34561 29365 34595
rect 29469 34561 29503 34595
rect 29561 34561 29595 34595
rect 29745 34561 29779 34595
rect 31401 34561 31435 34595
rect 32393 34561 32427 34595
rect 47593 34561 47627 34595
rect 21281 34493 21315 34527
rect 23673 34493 23707 34527
rect 23949 34493 23983 34527
rect 25605 34493 25639 34527
rect 29101 34493 29135 34527
rect 31585 34493 31619 34527
rect 32137 34493 32171 34527
rect 34345 34493 34379 34527
rect 34529 34493 34563 34527
rect 27169 34425 27203 34459
rect 47041 34425 47075 34459
rect 2053 34357 2087 34391
rect 24961 34357 24995 34391
rect 27905 34357 27939 34391
rect 28457 34357 28491 34391
rect 46397 34357 46431 34391
rect 47685 34357 47719 34391
rect 16313 34153 16347 34187
rect 18705 34153 18739 34187
rect 24777 34153 24811 34187
rect 25237 34153 25271 34187
rect 25973 34153 26007 34187
rect 26249 34153 26283 34187
rect 31401 34153 31435 34187
rect 34805 34153 34839 34187
rect 26985 34085 27019 34119
rect 1409 34017 1443 34051
rect 2789 34017 2823 34051
rect 24869 34017 24903 34051
rect 27537 34017 27571 34051
rect 46305 34017 46339 34051
rect 46489 34017 46523 34051
rect 48145 34017 48179 34051
rect 14933 33949 14967 33983
rect 16865 33949 16899 33983
rect 18337 33949 18371 33983
rect 21373 33949 21407 33983
rect 21649 33949 21683 33983
rect 25053 33949 25087 33983
rect 25881 33949 25915 33983
rect 26065 33949 26099 33983
rect 27445 33949 27479 33983
rect 28825 33949 28859 33983
rect 29561 33949 29595 33983
rect 31677 33949 31711 33983
rect 31769 33949 31803 33983
rect 31861 33949 31895 33983
rect 32045 33949 32079 33983
rect 32505 33949 32539 33983
rect 34713 33949 34747 33983
rect 1593 33881 1627 33915
rect 15200 33881 15234 33915
rect 16681 33881 16715 33915
rect 18521 33881 18555 33915
rect 23489 33881 23523 33915
rect 23673 33881 23707 33915
rect 24777 33881 24811 33915
rect 26801 33881 26835 33915
rect 28641 33881 28675 33915
rect 29806 33881 29840 33915
rect 32750 33881 32784 33915
rect 17049 33813 17083 33847
rect 23857 33813 23891 33847
rect 29009 33813 29043 33847
rect 30941 33813 30975 33847
rect 33885 33813 33919 33847
rect 2145 33609 2179 33643
rect 15485 33609 15519 33643
rect 18521 33609 18555 33643
rect 22385 33609 22419 33643
rect 28641 33609 28675 33643
rect 29009 33609 29043 33643
rect 32137 33609 32171 33643
rect 33425 33609 33459 33643
rect 46029 33609 46063 33643
rect 18429 33541 18463 33575
rect 22293 33541 22327 33575
rect 48145 33541 48179 33575
rect 2053 33473 2087 33507
rect 15761 33473 15795 33507
rect 15853 33473 15887 33507
rect 15945 33473 15979 33507
rect 16129 33473 16163 33507
rect 17509 33473 17543 33507
rect 17693 33473 17727 33507
rect 19625 33473 19659 33507
rect 23673 33473 23707 33507
rect 23765 33473 23799 33507
rect 23857 33473 23891 33507
rect 24041 33473 24075 33507
rect 25421 33473 25455 33507
rect 25513 33473 25547 33507
rect 25605 33473 25639 33507
rect 25789 33473 25823 33507
rect 27813 33473 27847 33507
rect 27997 33473 28031 33507
rect 28181 33473 28215 33507
rect 30113 33473 30147 33507
rect 30380 33473 30414 33507
rect 32413 33473 32447 33507
rect 32505 33473 32539 33507
rect 32597 33473 32631 33507
rect 32781 33473 32815 33507
rect 33333 33473 33367 33507
rect 45937 33473 45971 33507
rect 46581 33473 46615 33507
rect 47961 33473 47995 33507
rect 17233 33405 17267 33439
rect 29101 33405 29135 33439
rect 29193 33405 29227 33439
rect 19809 33337 19843 33371
rect 2881 33269 2915 33303
rect 17877 33269 17911 33303
rect 23397 33269 23431 33303
rect 25145 33269 25179 33303
rect 31493 33269 31527 33303
rect 46673 33269 46707 33303
rect 13461 33065 13495 33099
rect 23857 33065 23891 33099
rect 32597 33065 32631 33099
rect 17785 32997 17819 33031
rect 27169 32997 27203 33031
rect 28365 32997 28399 33031
rect 29561 32997 29595 33031
rect 13277 32929 13311 32963
rect 16405 32929 16439 32963
rect 21373 32929 21407 32963
rect 22937 32929 22971 32963
rect 24869 32929 24903 32963
rect 24961 32929 24995 32963
rect 30113 32929 30147 32963
rect 35173 32929 35207 32963
rect 37013 32929 37047 32963
rect 46305 32929 46339 32963
rect 46489 32929 46523 32963
rect 48053 32929 48087 32963
rect 2973 32861 3007 32895
rect 13185 32861 13219 32895
rect 14335 32861 14369 32895
rect 14470 32855 14504 32889
rect 14565 32861 14599 32895
rect 14749 32861 14783 32895
rect 18521 32861 18555 32895
rect 19901 32861 19935 32895
rect 19993 32861 20027 32895
rect 20085 32861 20119 32895
rect 20269 32861 20303 32895
rect 23489 32861 23523 32895
rect 25789 32861 25823 32895
rect 26045 32861 26079 32895
rect 27721 32861 27755 32895
rect 28641 32861 28675 32895
rect 28733 32861 28767 32895
rect 28825 32861 28859 32895
rect 29009 32861 29043 32895
rect 29929 32861 29963 32895
rect 32229 32861 32263 32895
rect 16672 32793 16706 32827
rect 18705 32793 18739 32827
rect 21189 32793 21223 32827
rect 22661 32793 22695 32827
rect 23673 32793 23707 32827
rect 27905 32793 27939 32827
rect 32413 32793 32447 32827
rect 35357 32793 35391 32827
rect 1869 32725 1903 32759
rect 3065 32725 3099 32759
rect 14105 32725 14139 32759
rect 19625 32725 19659 32759
rect 20729 32725 20763 32759
rect 21097 32725 21131 32759
rect 22293 32725 22327 32759
rect 22753 32725 22787 32759
rect 24409 32725 24443 32759
rect 24777 32725 24811 32759
rect 30021 32725 30055 32759
rect 12909 32521 12943 32555
rect 13645 32521 13679 32555
rect 16681 32521 16715 32555
rect 21005 32521 21039 32555
rect 25329 32521 25363 32555
rect 26341 32521 26375 32555
rect 14442 32453 14476 32487
rect 18153 32453 18187 32487
rect 30481 32453 30515 32487
rect 32229 32453 32263 32487
rect 1777 32385 1811 32419
rect 11785 32385 11819 32419
rect 13553 32385 13587 32419
rect 13737 32385 13771 32419
rect 16957 32385 16991 32419
rect 17046 32385 17080 32419
rect 17141 32388 17175 32422
rect 17325 32385 17359 32419
rect 17877 32385 17911 32419
rect 18061 32385 18095 32419
rect 19625 32385 19659 32419
rect 19892 32385 19926 32419
rect 21833 32385 21867 32419
rect 22089 32385 22123 32419
rect 23949 32385 23983 32419
rect 24205 32385 24239 32419
rect 25881 32385 25915 32419
rect 26157 32385 26191 32419
rect 27721 32385 27755 32419
rect 28365 32385 28399 32419
rect 28549 32385 28583 32419
rect 29561 32385 29595 32419
rect 32413 32385 32447 32419
rect 1961 32317 1995 32351
rect 2789 32317 2823 32351
rect 11529 32317 11563 32351
rect 14197 32317 14231 32351
rect 26065 32317 26099 32351
rect 29653 32317 29687 32351
rect 29837 32317 29871 32351
rect 27905 32249 27939 32283
rect 29193 32249 29227 32283
rect 30665 32249 30699 32283
rect 15577 32181 15611 32215
rect 23213 32181 23247 32215
rect 25881 32181 25915 32215
rect 28733 32181 28767 32215
rect 32597 32181 32631 32215
rect 10885 31977 10919 32011
rect 21925 31977 21959 32011
rect 31769 31977 31803 32011
rect 33885 31977 33919 32011
rect 35357 31977 35391 32011
rect 13553 31909 13587 31943
rect 27629 31909 27663 31943
rect 1409 31841 1443 31875
rect 1593 31841 1627 31875
rect 3893 31841 3927 31875
rect 10149 31841 10183 31875
rect 14105 31841 14139 31875
rect 14381 31841 14415 31875
rect 26157 31841 26191 31875
rect 28549 31841 28583 31875
rect 28733 31841 28767 31875
rect 30389 31841 30423 31875
rect 47869 31841 47903 31875
rect 3249 31773 3283 31807
rect 3801 31773 3835 31807
rect 10057 31773 10091 31807
rect 11161 31773 11195 31807
rect 11250 31773 11284 31807
rect 11345 31773 11379 31807
rect 11529 31773 11563 31807
rect 12173 31773 12207 31807
rect 17049 31773 17083 31807
rect 17233 31773 17267 31807
rect 17693 31773 17727 31807
rect 17877 31773 17911 31807
rect 18061 31773 18095 31807
rect 20637 31773 20671 31807
rect 20913 31773 20947 31807
rect 22155 31773 22189 31807
rect 22274 31770 22308 31804
rect 22374 31767 22408 31801
rect 22569 31773 22603 31807
rect 26433 31773 26467 31807
rect 26525 31773 26559 31807
rect 26638 31773 26672 31807
rect 26801 31773 26835 31807
rect 32505 31773 32539 31807
rect 35265 31773 35299 31807
rect 47501 31773 47535 31807
rect 12440 31705 12474 31739
rect 27261 31705 27295 31739
rect 27445 31705 27479 31739
rect 29561 31705 29595 31739
rect 29745 31705 29779 31739
rect 30634 31705 30668 31739
rect 32750 31705 32784 31739
rect 10425 31637 10459 31671
rect 28089 31637 28123 31671
rect 28457 31637 28491 31671
rect 29929 31637 29963 31671
rect 13093 31433 13127 31467
rect 13461 31433 13495 31467
rect 13553 31433 13587 31467
rect 22293 31433 22327 31467
rect 24317 31433 24351 31467
rect 25237 31433 25271 31467
rect 28549 31433 28583 31467
rect 29745 31433 29779 31467
rect 32137 31433 32171 31467
rect 1501 31365 1535 31399
rect 2329 31365 2363 31399
rect 14657 31365 14691 31399
rect 20361 31365 20395 31399
rect 21925 31365 21959 31399
rect 23213 31365 23247 31399
rect 27077 31365 27111 31399
rect 13369 31297 13403 31331
rect 14289 31297 14323 31331
rect 14473 31297 14507 31331
rect 16937 31297 16971 31331
rect 19717 31297 19751 31331
rect 20545 31297 20579 31331
rect 22109 31297 22143 31331
rect 23029 31297 23063 31331
rect 24225 31297 24259 31331
rect 25145 31297 25179 31331
rect 25881 31297 25915 31331
rect 28917 31297 28951 31331
rect 30021 31297 30055 31331
rect 30113 31297 30147 31331
rect 30205 31297 30239 31331
rect 30389 31297 30423 31331
rect 32413 31297 32447 31331
rect 32505 31297 32539 31331
rect 32597 31297 32631 31331
rect 32781 31297 32815 31331
rect 47961 31297 47995 31331
rect 2145 31229 2179 31263
rect 3157 31229 3191 31263
rect 13829 31229 13863 31263
rect 16681 31229 16715 31263
rect 20729 31229 20763 31263
rect 29009 31229 29043 31263
rect 29101 31229 29135 31263
rect 48145 31229 48179 31263
rect 19901 31161 19935 31195
rect 1593 31093 1627 31127
rect 13737 31093 13771 31127
rect 18061 31093 18095 31127
rect 23397 31093 23431 31127
rect 25973 31093 26007 31127
rect 27169 31093 27203 31127
rect 2329 30889 2363 30923
rect 3065 30889 3099 30923
rect 10333 30889 10367 30923
rect 16865 30889 16899 30923
rect 24409 30889 24443 30923
rect 40969 30889 41003 30923
rect 15209 30821 15243 30855
rect 22201 30753 22235 30787
rect 24869 30753 24903 30787
rect 24961 30753 24995 30787
rect 2237 30685 2271 30719
rect 10241 30685 10275 30719
rect 10425 30685 10459 30719
rect 11161 30685 11195 30719
rect 11250 30685 11284 30719
rect 11345 30685 11379 30719
rect 11529 30685 11563 30719
rect 14105 30685 14139 30719
rect 14289 30685 14323 30719
rect 16681 30685 16715 30719
rect 17601 30685 17635 30719
rect 17785 30685 17819 30719
rect 20591 30685 20625 30719
rect 20726 30685 20760 30719
rect 20821 30685 20855 30719
rect 21005 30685 21039 30719
rect 22017 30685 22051 30719
rect 23121 30685 23155 30719
rect 23213 30685 23247 30719
rect 23305 30685 23339 30719
rect 23489 30685 23523 30719
rect 25881 30685 25915 30719
rect 25973 30685 26007 30719
rect 26065 30685 26099 30719
rect 26249 30685 26283 30719
rect 26985 30685 27019 30719
rect 29837 30685 29871 30719
rect 29929 30685 29963 30719
rect 30021 30685 30055 30719
rect 30205 30685 30239 30719
rect 31401 30685 31435 30719
rect 33241 30685 33275 30719
rect 33977 30685 34011 30719
rect 34713 30685 34747 30719
rect 40785 30685 40819 30719
rect 10885 30617 10919 30651
rect 15025 30617 15059 30651
rect 19349 30617 19383 30651
rect 27230 30617 27264 30651
rect 31585 30617 31619 30651
rect 34069 30617 34103 30651
rect 34897 30617 34931 30651
rect 36553 30617 36587 30651
rect 14473 30549 14507 30583
rect 17141 30549 17175 30583
rect 17693 30549 17727 30583
rect 19441 30549 19475 30583
rect 20361 30549 20395 30583
rect 21649 30549 21683 30583
rect 22109 30549 22143 30583
rect 22845 30549 22879 30583
rect 24777 30549 24811 30583
rect 25605 30549 25639 30583
rect 28365 30549 28399 30583
rect 29561 30549 29595 30583
rect 31769 30549 31803 30583
rect 33333 30549 33367 30583
rect 10977 30345 11011 30379
rect 21281 30345 21315 30379
rect 24961 30345 24995 30379
rect 25881 30345 25915 30379
rect 13461 30277 13495 30311
rect 14289 30277 14323 30311
rect 14657 30277 14691 30311
rect 15393 30277 15427 30311
rect 16681 30277 16715 30311
rect 20913 30277 20947 30311
rect 33609 30277 33643 30311
rect 2237 30209 2271 30243
rect 7757 30209 7791 30243
rect 8024 30209 8058 30243
rect 9597 30209 9631 30243
rect 9864 30209 9898 30243
rect 13369 30209 13403 30243
rect 13553 30209 13587 30243
rect 14473 30209 14507 30243
rect 14749 30209 14783 30243
rect 15209 30209 15243 30243
rect 15485 30209 15519 30243
rect 16865 30209 16899 30243
rect 16957 30209 16991 30243
rect 17509 30209 17543 30243
rect 18153 30209 18187 30243
rect 21097 30209 21131 30243
rect 22937 30209 22971 30243
rect 23193 30209 23227 30243
rect 24869 30209 24903 30243
rect 25513 30209 25547 30243
rect 25697 30209 25731 30243
rect 31197 30209 31231 30243
rect 31306 30215 31340 30249
rect 31422 30209 31456 30243
rect 31585 30209 31619 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 33425 30209 33459 30243
rect 11621 30141 11655 30175
rect 11897 30141 11931 30175
rect 13829 30141 13863 30175
rect 18429 30141 18463 30175
rect 32505 30141 32539 30175
rect 35265 30141 35299 30175
rect 13737 30073 13771 30107
rect 15301 30073 15335 30107
rect 16681 30073 16715 30107
rect 1777 30005 1811 30039
rect 2329 30005 2363 30039
rect 9137 30005 9171 30039
rect 13093 30005 13127 30039
rect 17601 30005 17635 30039
rect 19533 30005 19567 30039
rect 24317 30005 24351 30039
rect 30941 30005 30975 30039
rect 10333 29801 10367 29835
rect 14105 29801 14139 29835
rect 18245 29801 18279 29835
rect 27629 29801 27663 29835
rect 33149 29801 33183 29835
rect 14565 29733 14599 29767
rect 1409 29665 1443 29699
rect 1593 29665 1627 29699
rect 2789 29665 2823 29699
rect 10977 29665 11011 29699
rect 11805 29665 11839 29699
rect 14197 29665 14231 29699
rect 17785 29665 17819 29699
rect 17877 29665 17911 29699
rect 28089 29665 28123 29699
rect 28181 29665 28215 29699
rect 31769 29665 31803 29699
rect 35541 29665 35575 29699
rect 47593 29665 47627 29699
rect 9505 29597 9539 29631
rect 10609 29597 10643 29631
rect 11069 29597 11103 29631
rect 11529 29597 11563 29631
rect 14381 29597 14415 29631
rect 15209 29597 15243 29631
rect 15393 29597 15427 29631
rect 17509 29597 17543 29631
rect 17697 29597 17731 29631
rect 18061 29597 18095 29631
rect 20729 29597 20763 29631
rect 20985 29597 21019 29631
rect 25789 29597 25823 29631
rect 30941 29597 30975 29631
rect 31033 29597 31067 29631
rect 31125 29597 31159 29631
rect 31309 29597 31343 29631
rect 32025 29597 32059 29631
rect 33609 29597 33643 29631
rect 34713 29597 34747 29631
rect 47317 29597 47351 29631
rect 9689 29529 9723 29563
rect 9873 29529 9907 29563
rect 10701 29529 10735 29563
rect 14105 29529 14139 29563
rect 15853 29529 15887 29563
rect 16037 29529 16071 29563
rect 19717 29529 19751 29563
rect 26034 29529 26068 29563
rect 35725 29529 35759 29563
rect 37381 29529 37415 29563
rect 10793 29461 10827 29495
rect 15301 29461 15335 29495
rect 16221 29461 16255 29495
rect 19809 29461 19843 29495
rect 22109 29461 22143 29495
rect 27169 29461 27203 29495
rect 27997 29461 28031 29495
rect 30665 29461 30699 29495
rect 33701 29461 33735 29495
rect 34805 29461 34839 29495
rect 9965 29257 9999 29291
rect 10885 29257 10919 29291
rect 11713 29257 11747 29291
rect 14749 29257 14783 29291
rect 30021 29257 30055 29291
rect 33609 29257 33643 29291
rect 37381 29257 37415 29291
rect 10517 29189 10551 29223
rect 10733 29189 10767 29223
rect 12992 29189 13026 29223
rect 23581 29189 23615 29223
rect 32474 29189 32508 29223
rect 2329 29121 2363 29155
rect 2973 29121 3007 29155
rect 9873 29121 9907 29155
rect 10057 29121 10091 29155
rect 11529 29121 11563 29155
rect 11805 29121 11839 29155
rect 12725 29121 12759 29155
rect 14657 29121 14691 29155
rect 15761 29121 15795 29155
rect 15853 29121 15887 29155
rect 15945 29121 15979 29155
rect 16129 29121 16163 29155
rect 16681 29121 16715 29155
rect 16937 29121 16971 29155
rect 19073 29121 19107 29155
rect 19257 29121 19291 29155
rect 23397 29121 23431 29155
rect 25697 29121 25731 29155
rect 28641 29121 28675 29155
rect 28908 29121 28942 29155
rect 31125 29121 31159 29155
rect 31217 29121 31251 29155
rect 31309 29121 31343 29155
rect 31493 29121 31527 29155
rect 32229 29121 32263 29155
rect 34529 29121 34563 29155
rect 37289 29121 37323 29155
rect 47593 29121 47627 29155
rect 25237 29053 25271 29087
rect 25789 29053 25823 29087
rect 34713 29053 34747 29087
rect 36369 29053 36403 29087
rect 11529 28985 11563 29019
rect 14105 28985 14139 29019
rect 18061 28985 18095 29019
rect 1869 28917 1903 28951
rect 2421 28917 2455 28951
rect 3065 28917 3099 28951
rect 10701 28917 10735 28951
rect 15485 28917 15519 28951
rect 19441 28917 19475 28951
rect 30849 28917 30883 28951
rect 47041 28917 47075 28951
rect 47685 28917 47719 28951
rect 17325 28713 17359 28747
rect 17509 28713 17543 28747
rect 23765 28713 23799 28747
rect 24593 28713 24627 28747
rect 25513 28713 25547 28747
rect 34805 28713 34839 28747
rect 18061 28645 18095 28679
rect 1409 28577 1443 28611
rect 2789 28577 2823 28611
rect 11253 28577 11287 28611
rect 12541 28577 12575 28611
rect 14289 28577 14323 28611
rect 14473 28577 14507 28611
rect 15761 28577 15795 28611
rect 16037 28577 16071 28611
rect 17233 28577 17267 28611
rect 19441 28577 19475 28611
rect 25697 28577 25731 28611
rect 26433 28577 26467 28611
rect 29929 28577 29963 28611
rect 30205 28577 30239 28611
rect 31217 28577 31251 28611
rect 37197 28577 37231 28611
rect 46305 28577 46339 28611
rect 48145 28577 48179 28611
rect 8401 28509 8435 28543
rect 9229 28509 9263 28543
rect 9321 28509 9355 28543
rect 9413 28509 9447 28543
rect 9597 28509 9631 28543
rect 10885 28509 10919 28543
rect 11345 28509 11379 28543
rect 12081 28509 12115 28543
rect 12449 28509 12483 28543
rect 13001 28509 13035 28543
rect 14381 28509 14415 28543
rect 14565 28509 14599 28543
rect 17325 28509 17359 28543
rect 18291 28509 18325 28543
rect 18429 28509 18463 28543
rect 18521 28509 18555 28543
rect 18705 28509 18739 28543
rect 23581 28509 23615 28543
rect 24409 28509 24443 28543
rect 25421 28509 25455 28543
rect 26157 28509 26191 28543
rect 31473 28509 31507 28543
rect 33333 28509 33367 28543
rect 34713 28509 34747 28543
rect 35541 28509 35575 28543
rect 1593 28441 1627 28475
rect 8033 28441 8067 28475
rect 8217 28441 8251 28475
rect 10977 28441 11011 28475
rect 12173 28441 12207 28475
rect 17049 28441 17083 28475
rect 19708 28441 19742 28475
rect 27997 28441 28031 28475
rect 28181 28441 28215 28475
rect 33885 28441 33919 28475
rect 35725 28441 35759 28475
rect 46489 28441 46523 28475
rect 8953 28373 8987 28407
rect 10609 28373 10643 28407
rect 11069 28373 11103 28407
rect 11805 28373 11839 28407
rect 12265 28373 12299 28407
rect 13093 28373 13127 28407
rect 14105 28373 14139 28407
rect 20821 28373 20855 28407
rect 25697 28373 25731 28407
rect 28365 28373 28399 28407
rect 32597 28373 32631 28407
rect 13001 28169 13035 28203
rect 14381 28169 14415 28203
rect 17233 28169 17267 28203
rect 17969 28169 18003 28203
rect 23213 28169 23247 28203
rect 37381 28169 37415 28203
rect 2881 28101 2915 28135
rect 9864 28101 9898 28135
rect 14013 28101 14047 28135
rect 19318 28101 19352 28135
rect 24041 28101 24075 28135
rect 24593 28101 24627 28135
rect 24777 28101 24811 28135
rect 34713 28101 34747 28135
rect 7113 28033 7147 28067
rect 7380 28033 7414 28067
rect 9597 28033 9631 28067
rect 12909 28033 12943 28067
rect 13093 28033 13127 28067
rect 14197 28033 14231 28067
rect 15117 28033 15151 28067
rect 17141 28033 17175 28067
rect 18225 28033 18259 28067
rect 18334 28033 18368 28067
rect 18429 28033 18463 28067
rect 18613 28033 18647 28067
rect 22477 28033 22511 28067
rect 23121 28033 23155 28067
rect 23857 28033 23891 28067
rect 25513 28033 25547 28067
rect 25605 28033 25639 28067
rect 25697 28033 25731 28067
rect 25881 28033 25915 28067
rect 27583 28033 27617 28067
rect 27721 28033 27755 28067
rect 27818 28033 27852 28067
rect 27997 28033 28031 28067
rect 29285 28033 29319 28067
rect 29377 28033 29411 28067
rect 29469 28033 29503 28067
rect 29653 28033 29687 28067
rect 30573 28033 30607 28067
rect 32781 28033 32815 28067
rect 34529 28033 34563 28067
rect 37289 28033 37323 28067
rect 47869 28033 47903 28067
rect 2697 27965 2731 27999
rect 4169 27965 4203 27999
rect 11529 27965 11563 27999
rect 11805 27965 11839 27999
rect 14841 27965 14875 27999
rect 19073 27965 19107 27999
rect 30941 27965 30975 27999
rect 33241 27965 33275 27999
rect 36369 27965 36403 27999
rect 10977 27897 11011 27931
rect 8493 27829 8527 27863
rect 20453 27829 20487 27863
rect 22569 27829 22603 27863
rect 25237 27829 25271 27863
rect 27353 27829 27387 27863
rect 29009 27829 29043 27863
rect 48053 27829 48087 27863
rect 17233 27625 17267 27659
rect 34897 27625 34931 27659
rect 8953 27557 8987 27591
rect 11161 27557 11195 27591
rect 16405 27557 16439 27591
rect 18061 27557 18095 27591
rect 21097 27557 21131 27591
rect 33885 27557 33919 27591
rect 11621 27489 11655 27523
rect 16589 27489 16623 27523
rect 25145 27489 25179 27523
rect 26801 27489 26835 27523
rect 29561 27489 29595 27523
rect 35633 27489 35667 27523
rect 37105 27489 37139 27523
rect 1593 27421 1627 27455
rect 2053 27421 2087 27455
rect 2881 27421 2915 27455
rect 6837 27421 6871 27455
rect 7104 27421 7138 27455
rect 9229 27421 9263 27455
rect 9321 27421 9355 27455
rect 9413 27421 9447 27455
rect 9597 27421 9631 27455
rect 10149 27421 10183 27455
rect 10333 27421 10367 27455
rect 11888 27421 11922 27455
rect 16313 27421 16347 27455
rect 17141 27421 17175 27455
rect 18317 27421 18351 27455
rect 18429 27421 18463 27455
rect 18542 27421 18576 27455
rect 18705 27421 18739 27455
rect 19717 27421 19751 27455
rect 21557 27421 21591 27455
rect 23397 27421 23431 27455
rect 24961 27421 24995 27455
rect 27261 27421 27295 27455
rect 27517 27421 27551 27455
rect 29817 27421 29851 27455
rect 31493 27421 31527 27455
rect 32413 27421 32447 27455
rect 34713 27421 34747 27455
rect 10793 27353 10827 27387
rect 10977 27353 11011 27387
rect 16589 27353 16623 27387
rect 19984 27353 20018 27387
rect 21802 27353 21836 27387
rect 31769 27353 31803 27387
rect 35817 27353 35851 27387
rect 2145 27285 2179 27319
rect 8217 27285 8251 27319
rect 10333 27285 10367 27319
rect 13001 27285 13035 27319
rect 22937 27285 22971 27319
rect 23581 27285 23615 27319
rect 28641 27285 28675 27319
rect 30941 27285 30975 27319
rect 8493 27081 8527 27115
rect 13553 27081 13587 27115
rect 13645 27081 13679 27115
rect 15577 27081 15611 27115
rect 19257 27081 19291 27115
rect 20085 27081 20119 27115
rect 29561 27081 29595 27115
rect 32505 27081 32539 27115
rect 35449 27081 35483 27115
rect 36185 27081 36219 27115
rect 37381 27081 37415 27115
rect 1961 27013 1995 27047
rect 17325 27013 17359 27047
rect 18889 27013 18923 27047
rect 19073 27013 19107 27047
rect 19901 27013 19935 27047
rect 22753 27013 22787 27047
rect 25320 27013 25354 27047
rect 27629 27013 27663 27047
rect 29193 27013 29227 27047
rect 32321 27013 32355 27047
rect 33149 27013 33183 27047
rect 1777 26945 1811 26979
rect 7113 26945 7147 26979
rect 8125 26945 8159 26979
rect 8309 26945 8343 26979
rect 13185 26945 13219 26979
rect 13461 26945 13495 26979
rect 13829 26945 13863 26979
rect 13921 26945 13955 26979
rect 15761 26945 15795 26979
rect 15945 26945 15979 26979
rect 17141 26945 17175 26979
rect 17417 26945 17451 26979
rect 19717 26945 19751 26979
rect 22569 26945 22603 26979
rect 25053 26945 25087 26979
rect 27445 26945 27479 26979
rect 28549 26945 28583 26979
rect 29377 26945 29411 26979
rect 30297 26945 30331 26979
rect 32137 26945 32171 26979
rect 32965 26945 32999 26979
rect 35265 26945 35299 26979
rect 36001 26945 36035 26979
rect 37289 26945 37323 26979
rect 37933 26945 37967 26979
rect 2789 26877 2823 26911
rect 14381 26877 14415 26911
rect 16037 26877 16071 26911
rect 23949 26877 23983 26911
rect 30665 26877 30699 26911
rect 34713 26877 34747 26911
rect 14749 26809 14783 26843
rect 7205 26741 7239 26775
rect 14841 26741 14875 26775
rect 17141 26741 17175 26775
rect 26433 26741 26467 26775
rect 28641 26741 28675 26775
rect 38025 26741 38059 26775
rect 16773 26537 16807 26571
rect 17233 26537 17267 26571
rect 18429 26537 18463 26571
rect 14749 26469 14783 26503
rect 17601 26469 17635 26503
rect 25145 26469 25179 26503
rect 1409 26401 1443 26435
rect 2789 26401 2823 26435
rect 6561 26401 6595 26435
rect 6745 26401 6779 26435
rect 7021 26401 7055 26435
rect 8953 26401 8987 26435
rect 10517 26401 10551 26435
rect 27813 26401 27847 26435
rect 28181 26401 28215 26435
rect 30849 26401 30883 26435
rect 32413 26401 32447 26435
rect 35541 26401 35575 26435
rect 35725 26401 35759 26435
rect 15393 26333 15427 26367
rect 17233 26333 17267 26367
rect 17417 26333 17451 26367
rect 18429 26333 18463 26367
rect 18705 26333 18739 26367
rect 19533 26333 19567 26367
rect 26157 26333 26191 26367
rect 27261 26333 27295 26367
rect 27445 26333 27479 26367
rect 28457 26333 28491 26367
rect 30205 26333 30239 26367
rect 31493 26333 31527 26367
rect 33517 26333 33551 26367
rect 34713 26333 34747 26367
rect 1593 26265 1627 26299
rect 9137 26265 9171 26299
rect 14565 26265 14599 26299
rect 15660 26265 15694 26299
rect 23673 26265 23707 26299
rect 24869 26265 24903 26299
rect 26525 26265 26559 26299
rect 34069 26265 34103 26299
rect 37381 26265 37415 26299
rect 47961 26265 47995 26299
rect 48145 26265 48179 26299
rect 18613 26197 18647 26231
rect 19717 26197 19751 26231
rect 23765 26197 23799 26231
rect 27353 26197 27387 26231
rect 34897 26197 34931 26231
rect 2329 25993 2363 26027
rect 8309 25993 8343 26027
rect 16681 25993 16715 26027
rect 17049 25993 17083 26027
rect 6377 25925 6411 25959
rect 26249 25925 26283 25959
rect 28273 25925 28307 25959
rect 29653 25925 29687 25959
rect 34713 25925 34747 25959
rect 1593 25857 1627 25891
rect 2237 25857 2271 25891
rect 6653 25857 6687 25891
rect 8217 25857 8251 25891
rect 9321 25857 9355 25891
rect 11713 25857 11747 25891
rect 13093 25857 13127 25891
rect 13277 25857 13311 25891
rect 14197 25857 14231 25891
rect 16865 25857 16899 25891
rect 17141 25857 17175 25891
rect 18512 25857 18546 25891
rect 20269 25857 20303 25891
rect 20453 25857 20487 25891
rect 20545 25857 20579 25891
rect 23489 25857 23523 25891
rect 23765 25857 23799 25891
rect 24593 25857 24627 25891
rect 25789 25857 25823 25891
rect 27077 25857 27111 25891
rect 27905 25857 27939 25891
rect 29469 25857 29503 25891
rect 32137 25857 32171 25891
rect 35173 25857 35207 25891
rect 6469 25789 6503 25823
rect 9597 25789 9631 25823
rect 11621 25789 11655 25823
rect 14289 25789 14323 25823
rect 18245 25789 18279 25823
rect 20085 25789 20119 25823
rect 23581 25789 23615 25823
rect 25145 25789 25179 25823
rect 31033 25789 31067 25823
rect 32873 25789 32907 25823
rect 33057 25789 33091 25823
rect 35817 25789 35851 25823
rect 1409 25721 1443 25755
rect 6377 25653 6411 25687
rect 6837 25653 6871 25687
rect 7297 25653 7331 25687
rect 11989 25653 12023 25687
rect 13185 25653 13219 25687
rect 19625 25653 19659 25687
rect 23489 25653 23523 25687
rect 23949 25653 23983 25687
rect 27261 25653 27295 25687
rect 32321 25653 32355 25687
rect 23213 25449 23247 25483
rect 23581 25449 23615 25483
rect 25513 25449 25547 25483
rect 11805 25381 11839 25415
rect 12081 25381 12115 25415
rect 24777 25381 24811 25415
rect 48053 25381 48087 25415
rect 9229 25313 9263 25347
rect 9689 25313 9723 25347
rect 10333 25313 10367 25347
rect 12173 25313 12207 25347
rect 13277 25313 13311 25347
rect 16221 25313 16255 25347
rect 20545 25313 20579 25347
rect 23213 25313 23247 25347
rect 8033 25245 8067 25279
rect 8125 25245 8159 25279
rect 8217 25245 8251 25279
rect 9597 25245 9631 25279
rect 10517 25245 10551 25279
rect 10609 25245 10643 25279
rect 10793 25245 10827 25279
rect 10885 25245 10919 25279
rect 11989 25245 12023 25279
rect 12265 25245 12299 25279
rect 13185 25245 13219 25279
rect 14105 25245 14139 25279
rect 14473 25245 14507 25279
rect 14565 25245 14599 25279
rect 16488 25245 16522 25279
rect 19257 25245 19291 25279
rect 19533 25245 19567 25279
rect 23397 25245 23431 25279
rect 24593 25245 24627 25279
rect 25329 25245 25363 25279
rect 26157 25245 26191 25279
rect 27997 25245 28031 25279
rect 29929 25245 29963 25279
rect 32321 25245 32355 25279
rect 33609 25245 33643 25279
rect 34713 25245 34747 25279
rect 47869 25245 47903 25279
rect 8401 25177 8435 25211
rect 9873 25177 9907 25211
rect 20812 25177 20846 25211
rect 23121 25177 23155 25211
rect 27261 25177 27295 25211
rect 28825 25177 28859 25211
rect 32965 25177 32999 25211
rect 13553 25109 13587 25143
rect 14381 25109 14415 25143
rect 17601 25109 17635 25143
rect 21925 25109 21959 25143
rect 31217 25109 31251 25143
rect 33793 25109 33827 25143
rect 34805 25109 34839 25143
rect 23489 24905 23523 24939
rect 8861 24837 8895 24871
rect 23949 24837 23983 24871
rect 24133 24837 24167 24871
rect 32229 24837 32263 24871
rect 7573 24769 7607 24803
rect 7757 24769 7791 24803
rect 8401 24769 8435 24803
rect 8585 24769 8619 24803
rect 9577 24769 9611 24803
rect 9670 24769 9704 24803
rect 9781 24772 9815 24806
rect 9965 24769 9999 24803
rect 10609 24769 10643 24803
rect 13461 24769 13495 24803
rect 18981 24769 19015 24803
rect 19165 24769 19199 24803
rect 19349 24769 19383 24803
rect 20683 24769 20717 24803
rect 20802 24775 20836 24809
rect 20913 24769 20947 24803
rect 21097 24769 21131 24803
rect 23018 24769 23052 24803
rect 23305 24769 23339 24803
rect 24961 24769 24995 24803
rect 25697 24769 25731 24803
rect 25881 24769 25915 24803
rect 27077 24769 27111 24803
rect 28089 24769 28123 24803
rect 28917 24769 28951 24803
rect 30757 24769 30791 24803
rect 32137 24769 32171 24803
rect 38025 24769 38059 24803
rect 38301 24769 38335 24803
rect 47593 24769 47627 24803
rect 7941 24701 7975 24735
rect 8769 24701 8803 24735
rect 10517 24701 10551 24735
rect 10977 24701 11011 24735
rect 13737 24701 13771 24735
rect 22753 24701 22787 24735
rect 23213 24701 23247 24735
rect 29285 24701 29319 24735
rect 30941 24701 30975 24735
rect 32781 24701 32815 24735
rect 32965 24701 32999 24735
rect 34437 24701 34471 24735
rect 38117 24701 38151 24735
rect 40049 24701 40083 24735
rect 40233 24701 40267 24735
rect 41245 24701 41279 24735
rect 20453 24633 20487 24667
rect 24317 24633 24351 24667
rect 8677 24565 8711 24599
rect 9321 24565 9355 24599
rect 13553 24565 13587 24599
rect 13645 24565 13679 24599
rect 23029 24565 23063 24599
rect 24133 24565 24167 24599
rect 25053 24565 25087 24599
rect 25973 24565 26007 24599
rect 27169 24565 27203 24599
rect 28181 24565 28215 24599
rect 38117 24565 38151 24599
rect 38485 24565 38519 24599
rect 47041 24565 47075 24599
rect 47685 24565 47719 24599
rect 9137 24361 9171 24395
rect 12909 24361 12943 24395
rect 22937 24361 22971 24395
rect 24409 24361 24443 24395
rect 40233 24361 40267 24395
rect 9965 24225 9999 24259
rect 24501 24225 24535 24259
rect 34713 24225 34747 24259
rect 34897 24225 34931 24259
rect 36553 24225 36587 24259
rect 46305 24225 46339 24259
rect 46489 24225 46523 24259
rect 48145 24225 48179 24259
rect 1409 24157 1443 24191
rect 9045 24157 9079 24191
rect 9229 24157 9263 24191
rect 9689 24157 9723 24191
rect 19717 24157 19751 24191
rect 24409 24157 24443 24191
rect 24685 24157 24719 24191
rect 25789 24157 25823 24191
rect 27629 24157 27663 24191
rect 29653 24157 29687 24191
rect 30757 24157 30791 24191
rect 31401 24157 31435 24191
rect 33241 24157 33275 24191
rect 33701 24157 33735 24191
rect 40141 24157 40175 24191
rect 12725 24089 12759 24123
rect 16405 24089 16439 24123
rect 16589 24089 16623 24123
rect 19984 24089 20018 24123
rect 21649 24089 21683 24123
rect 26034 24089 26068 24123
rect 27896 24089 27930 24123
rect 30021 24089 30055 24123
rect 30849 24089 30883 24123
rect 31585 24089 31619 24123
rect 1593 24021 1627 24055
rect 12925 24021 12959 24055
rect 13093 24021 13127 24055
rect 16773 24021 16807 24055
rect 21097 24021 21131 24055
rect 24869 24021 24903 24055
rect 27169 24021 27203 24055
rect 29009 24021 29043 24055
rect 33793 24021 33827 24055
rect 12725 23817 12759 23851
rect 20361 23817 20395 23851
rect 23121 23817 23155 23851
rect 25789 23817 25823 23851
rect 27353 23817 27387 23851
rect 27905 23817 27939 23851
rect 31585 23817 31619 23851
rect 32689 23817 32723 23851
rect 48053 23817 48087 23851
rect 14289 23749 14323 23783
rect 19257 23749 19291 23783
rect 19441 23749 19475 23783
rect 19625 23749 19659 23783
rect 47961 23749 47995 23783
rect 7389 23681 7423 23715
rect 9689 23681 9723 23715
rect 9781 23681 9815 23715
rect 11713 23681 11747 23715
rect 12541 23681 12575 23715
rect 12817 23681 12851 23715
rect 13461 23681 13495 23715
rect 14565 23681 14599 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 17141 23681 17175 23715
rect 17325 23681 17359 23715
rect 18107 23681 18141 23715
rect 18226 23681 18260 23715
rect 18337 23681 18371 23715
rect 18521 23681 18555 23715
rect 20637 23681 20671 23715
rect 20726 23681 20760 23715
rect 20826 23681 20860 23715
rect 21005 23681 21039 23715
rect 23213 23681 23247 23715
rect 23305 23681 23339 23715
rect 24133 23681 24167 23715
rect 24225 23681 24259 23715
rect 24685 23681 24719 23715
rect 26019 23681 26053 23715
rect 26154 23681 26188 23715
rect 26249 23681 26283 23715
rect 26433 23681 26467 23715
rect 26985 23681 27019 23715
rect 27169 23681 27203 23715
rect 28181 23681 28215 23715
rect 28273 23681 28307 23715
rect 28365 23681 28399 23715
rect 28549 23681 28583 23715
rect 29377 23681 29411 23715
rect 29561 23681 29595 23715
rect 30472 23681 30506 23715
rect 32597 23681 32631 23715
rect 7573 23613 7607 23647
rect 9137 23613 9171 23647
rect 9965 23613 9999 23647
rect 11621 23613 11655 23647
rect 13553 23613 13587 23647
rect 14381 23613 14415 23647
rect 24593 23613 24627 23647
rect 30205 23613 30239 23647
rect 33241 23613 33275 23647
rect 33425 23613 33459 23647
rect 33793 23613 33827 23647
rect 12081 23545 12115 23579
rect 13829 23545 13863 23579
rect 22937 23545 22971 23579
rect 2053 23477 2087 23511
rect 9873 23477 9907 23511
rect 12541 23477 12575 23511
rect 14473 23477 14507 23511
rect 14749 23477 14783 23511
rect 16681 23477 16715 23511
rect 17877 23477 17911 23511
rect 23489 23477 23523 23511
rect 29745 23477 29779 23511
rect 7849 23273 7883 23307
rect 9505 23273 9539 23307
rect 9689 23273 9723 23307
rect 10701 23273 10735 23307
rect 12541 23273 12575 23307
rect 13001 23273 13035 23307
rect 14289 23273 14323 23307
rect 14473 23273 14507 23307
rect 24409 23273 24443 23307
rect 28825 23273 28859 23307
rect 29929 23273 29963 23307
rect 16957 23205 16991 23239
rect 18061 23205 18095 23239
rect 20545 23205 20579 23239
rect 24869 23205 24903 23239
rect 1409 23137 1443 23171
rect 2789 23137 2823 23171
rect 10425 23137 10459 23171
rect 12633 23137 12667 23171
rect 24501 23137 24535 23171
rect 7757 23069 7791 23103
rect 9321 23069 9355 23103
rect 9505 23069 9539 23103
rect 10333 23069 10367 23103
rect 12541 23069 12575 23103
rect 12817 23069 12851 23103
rect 15577 23069 15611 23103
rect 15844 23069 15878 23103
rect 17877 23069 17911 23103
rect 20177 23069 20211 23103
rect 23673 23069 23707 23103
rect 23857 23069 23891 23103
rect 24685 23069 24719 23103
rect 25329 23069 25363 23103
rect 28641 23069 28675 23103
rect 30205 23069 30239 23103
rect 30294 23069 30328 23103
rect 30389 23069 30423 23103
rect 30573 23069 30607 23103
rect 31033 23069 31067 23103
rect 1593 23001 1627 23035
rect 14131 23001 14165 23035
rect 14321 23001 14355 23035
rect 17693 23001 17727 23035
rect 20361 23001 20395 23035
rect 21097 23001 21131 23035
rect 23765 23001 23799 23035
rect 24409 23001 24443 23035
rect 28457 23001 28491 23035
rect 21189 22933 21223 22967
rect 25513 22933 25547 22967
rect 31125 22933 31159 22967
rect 2605 22729 2639 22763
rect 31585 22729 31619 22763
rect 12817 22661 12851 22695
rect 13645 22661 13679 22695
rect 14289 22661 14323 22695
rect 16957 22661 16991 22695
rect 17684 22661 17718 22695
rect 23857 22661 23891 22695
rect 26157 22661 26191 22695
rect 1869 22593 1903 22627
rect 2513 22593 2547 22627
rect 12725 22593 12759 22627
rect 12909 22593 12943 22627
rect 13369 22593 13403 22627
rect 14105 22593 14139 22627
rect 14381 22593 14415 22627
rect 16773 22593 16807 22627
rect 19533 22593 19567 22627
rect 20545 22593 20579 22627
rect 20729 22593 20763 22627
rect 21833 22593 21867 22627
rect 22100 22593 22134 22627
rect 23765 22593 23799 22627
rect 24869 22593 24903 22627
rect 25145 22593 25179 22627
rect 26985 22593 27019 22627
rect 27261 22593 27295 22627
rect 29331 22593 29365 22627
rect 29469 22593 29503 22627
rect 29561 22593 29595 22627
rect 29745 22593 29779 22627
rect 30205 22593 30239 22627
rect 30461 22593 30495 22627
rect 34069 22593 34103 22627
rect 34161 22593 34195 22627
rect 34253 22593 34287 22627
rect 34437 22593 34471 22627
rect 48145 22593 48179 22627
rect 13461 22525 13495 22559
rect 13645 22525 13679 22559
rect 17417 22525 17451 22559
rect 19257 22525 19291 22559
rect 25053 22525 25087 22559
rect 14105 22457 14139 22491
rect 18797 22457 18831 22491
rect 29101 22457 29135 22491
rect 1961 22389 1995 22423
rect 20913 22389 20947 22423
rect 23213 22389 23247 22423
rect 25145 22389 25179 22423
rect 25329 22389 25363 22423
rect 26249 22389 26283 22423
rect 33793 22389 33827 22423
rect 47961 22389 47995 22423
rect 14289 22185 14323 22219
rect 23673 22185 23707 22219
rect 24409 22185 24443 22219
rect 24869 22185 24903 22219
rect 47869 22185 47903 22219
rect 14473 22117 14507 22151
rect 10885 22049 10919 22083
rect 29745 22049 29779 22083
rect 33057 22049 33091 22083
rect 47409 22049 47443 22083
rect 9137 21981 9171 22015
rect 10241 21981 10275 22015
rect 14105 21981 14139 22015
rect 14289 21981 14323 22015
rect 18291 21981 18325 22015
rect 18429 21981 18463 22015
rect 18521 21981 18555 22015
rect 18705 21981 18739 22015
rect 19257 21981 19291 22015
rect 21419 21981 21453 22015
rect 21554 21981 21588 22015
rect 21649 21981 21683 22015
rect 21833 21981 21867 22015
rect 23673 21981 23707 22015
rect 23857 21981 23891 22015
rect 24593 21981 24627 22015
rect 24685 21981 24719 22015
rect 25605 21981 25639 22015
rect 27629 21981 27663 22015
rect 29561 21981 29595 22015
rect 33793 21981 33827 22015
rect 33885 21981 33919 22015
rect 33977 21981 34011 22015
rect 34161 21981 34195 22015
rect 34713 21981 34747 22015
rect 47501 21981 47535 22015
rect 47869 21981 47903 22015
rect 8953 21913 8987 21947
rect 11069 21913 11103 21947
rect 12725 21913 12759 21947
rect 18061 21913 18095 21947
rect 19502 21913 19536 21947
rect 21189 21913 21223 21947
rect 24409 21913 24443 21947
rect 25850 21913 25884 21947
rect 27896 21913 27930 21947
rect 31401 21913 31435 21947
rect 32689 21913 32723 21947
rect 32873 21913 32907 21947
rect 34958 21913 34992 21947
rect 9321 21845 9355 21879
rect 10333 21845 10367 21879
rect 20637 21845 20671 21879
rect 26985 21845 27019 21879
rect 29009 21845 29043 21879
rect 33517 21845 33551 21879
rect 36093 21845 36127 21879
rect 48053 21845 48087 21879
rect 8861 21641 8895 21675
rect 11621 21641 11655 21675
rect 13461 21641 13495 21675
rect 19349 21641 19383 21675
rect 28273 21641 28307 21675
rect 30573 21641 30607 21675
rect 7748 21573 7782 21607
rect 9321 21573 9355 21607
rect 19165 21573 19199 21607
rect 20729 21573 20763 21607
rect 26985 21573 27019 21607
rect 29377 21573 29411 21607
rect 29561 21573 29595 21607
rect 47961 21573 47995 21607
rect 9597 21505 9631 21539
rect 9689 21505 9723 21539
rect 9781 21505 9815 21539
rect 9965 21505 9999 21539
rect 11529 21505 11563 21539
rect 13001 21505 13035 21539
rect 13277 21505 13311 21539
rect 17141 21505 17175 21539
rect 17877 21505 17911 21539
rect 18981 21505 19015 21539
rect 19993 21505 20027 21539
rect 22365 21505 22399 21539
rect 23949 21505 23983 21539
rect 25651 21505 25685 21539
rect 25789 21505 25823 21539
rect 25881 21505 25915 21539
rect 26065 21505 26099 21539
rect 27169 21505 27203 21539
rect 28503 21505 28537 21539
rect 28641 21505 28675 21539
rect 28733 21505 28767 21539
rect 28917 21505 28951 21539
rect 30205 21505 30239 21539
rect 30389 21505 30423 21539
rect 33793 21505 33827 21539
rect 34049 21505 34083 21539
rect 7481 21437 7515 21471
rect 13185 21437 13219 21471
rect 14013 21437 14047 21471
rect 14289 21437 14323 21471
rect 22109 21437 22143 21471
rect 25421 21437 25455 21471
rect 27353 21437 27387 21471
rect 29745 21437 29779 21471
rect 17325 21369 17359 21403
rect 20913 21369 20947 21403
rect 13277 21301 13311 21335
rect 17969 21301 18003 21335
rect 19809 21301 19843 21335
rect 23489 21301 23523 21335
rect 24179 21301 24213 21335
rect 35173 21301 35207 21335
rect 48053 21301 48087 21335
rect 33977 21097 34011 21131
rect 15669 21029 15703 21063
rect 20913 21029 20947 21063
rect 21373 21029 21407 21063
rect 6929 20961 6963 20995
rect 10609 20961 10643 20995
rect 11069 20961 11103 20995
rect 24777 20961 24811 20995
rect 26893 20961 26927 20995
rect 6285 20893 6319 20927
rect 9183 20893 9217 20927
rect 9318 20890 9352 20924
rect 9413 20893 9447 20927
rect 9597 20893 9631 20927
rect 10425 20893 10459 20927
rect 14289 20893 14323 20927
rect 16129 20893 16163 20927
rect 19717 20893 19751 20927
rect 20729 20893 20763 20927
rect 21649 20893 21683 20927
rect 21754 20887 21788 20921
rect 21854 20893 21888 20927
rect 22017 20893 22051 20927
rect 24409 20893 24443 20927
rect 26249 20893 26283 20927
rect 31539 20893 31573 20927
rect 31677 20893 31711 20927
rect 31790 20890 31824 20924
rect 31953 20893 31987 20927
rect 32597 20893 32631 20927
rect 33609 20893 33643 20927
rect 33793 20893 33827 20927
rect 6469 20825 6503 20859
rect 14556 20825 14590 20859
rect 16396 20825 16430 20859
rect 22569 20825 22603 20859
rect 23673 20825 23707 20859
rect 24593 20825 24627 20859
rect 26341 20825 26375 20859
rect 27077 20825 27111 20859
rect 28733 20825 28767 20859
rect 32413 20825 32447 20859
rect 8953 20757 8987 20791
rect 17509 20757 17543 20791
rect 19809 20757 19843 20791
rect 22661 20757 22695 20791
rect 23765 20757 23799 20791
rect 31309 20757 31343 20791
rect 32781 20757 32815 20791
rect 6469 20553 6503 20587
rect 8769 20553 8803 20587
rect 9597 20553 9631 20587
rect 14473 20553 14507 20587
rect 16681 20553 16715 20587
rect 18245 20485 18279 20519
rect 27997 20485 28031 20519
rect 28181 20485 28215 20519
rect 6377 20417 6411 20451
rect 7389 20417 7423 20451
rect 7656 20417 7690 20451
rect 9229 20417 9263 20451
rect 9413 20417 9447 20451
rect 10609 20417 10643 20451
rect 10793 20417 10827 20451
rect 10977 20417 11011 20451
rect 12219 20417 12253 20451
rect 12357 20417 12391 20451
rect 12449 20417 12483 20451
rect 12633 20417 12667 20451
rect 13645 20417 13679 20451
rect 13737 20417 13771 20451
rect 13829 20417 13863 20451
rect 14013 20417 14047 20451
rect 14749 20417 14783 20451
rect 14838 20417 14872 20451
rect 14933 20417 14967 20451
rect 15117 20417 15151 20451
rect 15669 20417 15703 20451
rect 15853 20417 15887 20451
rect 16957 20417 16991 20451
rect 17049 20417 17083 20451
rect 17141 20417 17175 20451
rect 17325 20417 17359 20451
rect 18061 20417 18095 20451
rect 19625 20417 19659 20451
rect 20545 20417 20579 20451
rect 20637 20417 20671 20451
rect 20729 20417 20763 20451
rect 20913 20417 20947 20451
rect 23305 20417 23339 20451
rect 30205 20417 30239 20451
rect 30461 20417 30495 20451
rect 32137 20417 32171 20451
rect 32393 20417 32427 20451
rect 34253 20417 34287 20451
rect 34345 20417 34379 20451
rect 34437 20417 34471 20451
rect 34621 20417 34655 20451
rect 31585 20281 31619 20315
rect 33517 20281 33551 20315
rect 11989 20213 12023 20247
rect 13369 20213 13403 20247
rect 16037 20213 16071 20247
rect 17693 20213 17727 20247
rect 18429 20213 18463 20247
rect 19717 20213 19751 20247
rect 20269 20213 20303 20247
rect 23397 20213 23431 20247
rect 33977 20213 34011 20247
rect 11529 20009 11563 20043
rect 13553 20009 13587 20043
rect 14473 20009 14507 20043
rect 20637 19941 20671 19975
rect 25789 19941 25823 19975
rect 26525 19941 26559 19975
rect 34069 19941 34103 19975
rect 34713 19873 34747 19907
rect 46305 19873 46339 19907
rect 2053 19805 2087 19839
rect 10149 19805 10183 19839
rect 10416 19805 10450 19839
rect 12173 19805 12207 19839
rect 13185 19805 13219 19839
rect 14289 19805 14323 19839
rect 16957 19805 16991 19839
rect 17049 19805 17083 19839
rect 17162 19805 17196 19839
rect 17325 19805 17359 19839
rect 18291 19805 18325 19839
rect 18429 19805 18463 19839
rect 18521 19805 18555 19839
rect 18705 19805 18739 19839
rect 19257 19805 19291 19839
rect 21189 19805 21223 19839
rect 21456 19805 21490 19839
rect 24409 19805 24443 19839
rect 27997 19805 28031 19839
rect 29561 19805 29595 19839
rect 31585 19805 31619 19839
rect 32229 19805 32263 19839
rect 32413 19805 32447 19839
rect 33701 19805 33735 19839
rect 33885 19805 33919 19839
rect 34969 19805 35003 19839
rect 11989 19737 12023 19771
rect 13369 19737 13403 19771
rect 14105 19737 14139 19771
rect 18061 19737 18095 19771
rect 19502 19737 19536 19771
rect 24676 19737 24710 19771
rect 26341 19737 26375 19771
rect 27813 19737 27847 19771
rect 29806 19737 29840 19771
rect 31401 19737 31435 19771
rect 46489 19737 46523 19771
rect 48145 19737 48179 19771
rect 12357 19669 12391 19703
rect 16681 19669 16715 19703
rect 22569 19669 22603 19703
rect 30941 19669 30975 19703
rect 31769 19669 31803 19703
rect 32597 19669 32631 19703
rect 36093 19669 36127 19703
rect 14565 19465 14599 19499
rect 18153 19465 18187 19499
rect 26065 19465 26099 19499
rect 28641 19465 28675 19499
rect 30297 19465 30331 19499
rect 33609 19465 33643 19499
rect 46765 19465 46799 19499
rect 10793 19397 10827 19431
rect 16129 19397 16163 19431
rect 18889 19397 18923 19431
rect 22293 19397 22327 19431
rect 23213 19397 23247 19431
rect 1869 19329 1903 19363
rect 7757 19329 7791 19363
rect 12357 19329 12391 19363
rect 12462 19335 12496 19369
rect 12562 19329 12596 19363
rect 12725 19329 12759 19363
rect 13185 19329 13219 19363
rect 13452 19329 13486 19363
rect 15945 19329 15979 19363
rect 16773 19329 16807 19363
rect 17029 19329 17063 19363
rect 18705 19329 18739 19363
rect 19809 19329 19843 19363
rect 19993 19329 20027 19363
rect 23029 19329 23063 19363
rect 25329 19329 25363 19363
rect 26249 19329 26283 19363
rect 28917 19329 28951 19363
rect 29009 19329 29043 19363
rect 29101 19329 29135 19363
rect 29285 19329 29319 19363
rect 30527 19329 30561 19363
rect 30662 19335 30696 19369
rect 30757 19329 30791 19363
rect 30941 19329 30975 19363
rect 32229 19329 32263 19363
rect 32485 19329 32519 19363
rect 46673 19329 46707 19363
rect 2053 19261 2087 19295
rect 2789 19261 2823 19295
rect 7941 19261 7975 19295
rect 8217 19261 8251 19295
rect 10977 19261 11011 19295
rect 23949 19261 23983 19295
rect 25605 19261 25639 19295
rect 47777 19261 47811 19295
rect 20177 19193 20211 19227
rect 12081 19125 12115 19159
rect 22385 19125 22419 19159
rect 25421 19125 25455 19159
rect 25513 19125 25547 19159
rect 2329 18921 2363 18955
rect 8125 18921 8159 18955
rect 11805 18921 11839 18955
rect 17601 18921 17635 18955
rect 24777 18921 24811 18955
rect 26433 18921 26467 18955
rect 29009 18921 29043 18955
rect 30113 18921 30147 18955
rect 31585 18921 31619 18955
rect 12265 18785 12299 18819
rect 22753 18785 22787 18819
rect 25329 18785 25363 18819
rect 47317 18785 47351 18819
rect 47593 18785 47627 18819
rect 2237 18717 2271 18751
rect 7113 18717 7147 18751
rect 8033 18717 8067 18751
rect 9229 18717 9263 18751
rect 9321 18717 9355 18751
rect 9413 18717 9447 18751
rect 9597 18717 9631 18751
rect 10425 18717 10459 18751
rect 10692 18717 10726 18751
rect 12541 18717 12575 18751
rect 15761 18717 15795 18751
rect 16037 18717 16071 18751
rect 17233 18717 17267 18751
rect 17417 18717 17451 18751
rect 22477 18717 22511 18751
rect 22569 18717 22603 18751
rect 26157 18717 26191 18751
rect 26249 18717 26283 18751
rect 26525 18717 26559 18751
rect 28181 18717 28215 18751
rect 30021 18717 30055 18751
rect 31861 18717 31895 18751
rect 31953 18717 31987 18751
rect 32045 18717 32079 18751
rect 32229 18717 32263 18751
rect 25145 18649 25179 18683
rect 27997 18649 28031 18683
rect 28641 18649 28675 18683
rect 28825 18649 28859 18683
rect 7205 18581 7239 18615
rect 8953 18581 8987 18615
rect 22753 18581 22787 18615
rect 25237 18581 25271 18615
rect 25973 18581 26007 18615
rect 25145 18377 25179 18411
rect 25605 18377 25639 18411
rect 26065 18377 26099 18411
rect 6745 18309 6779 18343
rect 6837 18309 6871 18343
rect 8116 18309 8150 18343
rect 10609 18309 10643 18343
rect 10977 18309 11011 18343
rect 15669 18309 15703 18343
rect 16773 18309 16807 18343
rect 19165 18309 19199 18343
rect 2053 18241 2087 18275
rect 2697 18241 2731 18275
rect 10793 18241 10827 18275
rect 12035 18241 12069 18275
rect 12170 18244 12204 18278
rect 12265 18244 12299 18278
rect 12449 18241 12483 18275
rect 13691 18241 13725 18275
rect 13842 18241 13876 18275
rect 13942 18241 13976 18275
rect 14105 18241 14139 18275
rect 14657 18241 14691 18275
rect 15485 18241 15519 18275
rect 18245 18241 18279 18275
rect 18334 18241 18368 18275
rect 18450 18241 18484 18275
rect 18613 18241 18647 18275
rect 19349 18241 19383 18275
rect 21833 18241 21867 18275
rect 22100 18241 22134 18275
rect 23673 18241 23707 18275
rect 24777 18241 24811 18275
rect 24961 18241 24995 18275
rect 25973 18241 26007 18275
rect 27629 18241 27663 18275
rect 27896 18241 27930 18275
rect 7849 18173 7883 18207
rect 23765 18173 23799 18207
rect 26157 18173 26191 18207
rect 7297 18105 7331 18139
rect 1593 18037 1627 18071
rect 2145 18037 2179 18071
rect 2789 18037 2823 18071
rect 9229 18037 9263 18071
rect 11805 18037 11839 18071
rect 13461 18037 13495 18071
rect 14749 18037 14783 18071
rect 16865 18037 16899 18071
rect 17969 18037 18003 18071
rect 19533 18037 19567 18071
rect 23213 18037 23247 18071
rect 23857 18037 23891 18071
rect 24041 18037 24075 18071
rect 29009 18037 29043 18071
rect 7573 17833 7607 17867
rect 8401 17833 8435 17867
rect 12081 17833 12115 17867
rect 13553 17833 13587 17867
rect 18061 17833 18095 17867
rect 20637 17833 20671 17867
rect 24777 17833 24811 17867
rect 25697 17833 25731 17867
rect 29929 17833 29963 17867
rect 16589 17765 16623 17799
rect 17601 17765 17635 17799
rect 21925 17765 21959 17799
rect 22569 17765 22603 17799
rect 26065 17765 26099 17799
rect 27261 17765 27295 17799
rect 28549 17765 28583 17799
rect 1409 17697 1443 17731
rect 2789 17697 2823 17731
rect 15301 17697 15335 17731
rect 19257 17697 19291 17731
rect 21787 17697 21821 17731
rect 23213 17697 23247 17731
rect 27721 17697 27755 17731
rect 27813 17697 27847 17731
rect 28733 17697 28767 17731
rect 30021 17697 30055 17731
rect 7205 17629 7239 17663
rect 8217 17629 8251 17663
rect 9229 17629 9263 17663
rect 9321 17629 9355 17663
rect 9413 17629 9447 17663
rect 9597 17629 9631 17663
rect 10701 17629 10735 17663
rect 10968 17629 11002 17663
rect 13185 17629 13219 17663
rect 13369 17629 13403 17663
rect 14197 17629 14231 17663
rect 15025 17629 15059 17663
rect 16405 17629 16439 17663
rect 18337 17629 18371 17663
rect 18426 17629 18460 17663
rect 18521 17629 18555 17663
rect 18705 17629 18739 17663
rect 19513 17629 19547 17663
rect 21649 17629 21683 17663
rect 22109 17629 22143 17663
rect 23029 17629 23063 17663
rect 24501 17629 24535 17663
rect 24685 17629 24719 17663
rect 24777 17629 24811 17663
rect 25881 17629 25915 17663
rect 26157 17629 26191 17663
rect 27629 17629 27663 17663
rect 28457 17629 28491 17663
rect 29745 17629 29779 17663
rect 47685 17629 47719 17663
rect 1593 17561 1627 17595
rect 7389 17561 7423 17595
rect 8033 17561 8067 17595
rect 14381 17561 14415 17595
rect 17417 17561 17451 17595
rect 8953 17493 8987 17527
rect 14565 17493 14599 17527
rect 22109 17493 22143 17527
rect 22937 17493 22971 17527
rect 24961 17493 24995 17527
rect 28733 17493 28767 17527
rect 29561 17493 29595 17527
rect 9229 17289 9263 17323
rect 20269 17289 20303 17323
rect 22569 17289 22603 17323
rect 23489 17289 23523 17323
rect 25145 17289 25179 17323
rect 26341 17289 26375 17323
rect 30021 17289 30055 17323
rect 1593 17221 1627 17255
rect 24685 17221 24719 17255
rect 29101 17221 29135 17255
rect 3709 17153 3743 17187
rect 7849 17153 7883 17187
rect 8116 17153 8150 17187
rect 13452 17153 13486 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 15669 17153 15703 17187
rect 16773 17153 16807 17187
rect 16957 17153 16991 17187
rect 17417 17153 17451 17187
rect 17601 17153 17635 17187
rect 18061 17153 18095 17187
rect 18317 17153 18351 17187
rect 20177 17153 20211 17187
rect 21833 17153 21867 17187
rect 22937 17153 22971 17187
rect 23029 17153 23063 17187
rect 23213 17153 23247 17187
rect 23673 17153 23707 17187
rect 23765 17153 23799 17187
rect 24961 17153 24995 17187
rect 26157 17153 26191 17187
rect 28917 17153 28951 17187
rect 29193 17153 29227 17187
rect 32137 17153 32171 17187
rect 32404 17153 32438 17187
rect 47593 17153 47627 17187
rect 1409 17085 1443 17119
rect 2789 17085 2823 17119
rect 3893 17085 3927 17119
rect 4169 17085 4203 17119
rect 13185 17085 13219 17119
rect 15025 17085 15059 17119
rect 22109 17085 22143 17119
rect 23857 17085 23891 17119
rect 23949 17085 23983 17119
rect 24869 17085 24903 17119
rect 27445 17085 27479 17119
rect 27721 17085 27755 17119
rect 30113 17085 30147 17119
rect 30297 17085 30331 17119
rect 14565 17017 14599 17051
rect 19441 17017 19475 17051
rect 22017 17017 22051 17051
rect 28733 17017 28767 17051
rect 16865 16949 16899 16983
rect 17509 16949 17543 16983
rect 21925 16949 21959 16983
rect 24317 16949 24351 16983
rect 24685 16949 24719 16983
rect 29653 16949 29687 16983
rect 33517 16949 33551 16983
rect 47041 16949 47075 16983
rect 47685 16949 47719 16983
rect 2697 16745 2731 16779
rect 3893 16745 3927 16779
rect 17417 16745 17451 16779
rect 19625 16745 19659 16779
rect 23673 16745 23707 16779
rect 25329 16745 25363 16779
rect 28273 16745 28307 16779
rect 33517 16745 33551 16779
rect 2053 16677 2087 16711
rect 29009 16677 29043 16711
rect 30389 16677 30423 16711
rect 10977 16609 11011 16643
rect 11437 16609 11471 16643
rect 15393 16609 15427 16643
rect 22661 16609 22695 16643
rect 22845 16609 22879 16643
rect 23489 16609 23523 16643
rect 25881 16609 25915 16643
rect 27905 16609 27939 16643
rect 30941 16609 30975 16643
rect 33057 16609 33091 16643
rect 33149 16609 33183 16643
rect 46305 16609 46339 16643
rect 48145 16609 48179 16643
rect 1869 16541 1903 16575
rect 3801 16541 3835 16575
rect 14565 16541 14599 16575
rect 14657 16541 14691 16575
rect 14754 16541 14788 16575
rect 14933 16541 14967 16575
rect 17325 16541 17359 16575
rect 18521 16541 18555 16575
rect 20637 16541 20671 16575
rect 21281 16541 21315 16575
rect 23397 16541 23431 16575
rect 23673 16541 23707 16575
rect 26157 16541 26191 16575
rect 27537 16541 27571 16575
rect 27721 16541 27755 16575
rect 27813 16541 27847 16575
rect 28089 16541 28123 16575
rect 29837 16541 29871 16575
rect 30021 16541 30055 16575
rect 30205 16541 30239 16575
rect 32781 16541 32815 16575
rect 32965 16541 32999 16575
rect 33333 16541 33367 16575
rect 11161 16473 11195 16507
rect 15638 16473 15672 16507
rect 18705 16473 18739 16507
rect 19257 16473 19291 16507
rect 19441 16473 19475 16507
rect 22569 16473 22603 16507
rect 25053 16473 25087 16507
rect 28825 16473 28859 16507
rect 30113 16473 30147 16507
rect 31186 16473 31220 16507
rect 46489 16473 46523 16507
rect 14289 16405 14323 16439
rect 16773 16405 16807 16439
rect 22201 16405 22235 16439
rect 23857 16405 23891 16439
rect 32321 16405 32355 16439
rect 11621 16201 11655 16235
rect 17509 16201 17543 16235
rect 18705 16201 18739 16235
rect 21925 16201 21959 16235
rect 29009 16201 29043 16235
rect 30481 16201 30515 16235
rect 24041 16133 24075 16167
rect 24593 16133 24627 16167
rect 24777 16133 24811 16167
rect 25421 16133 25455 16167
rect 27997 16133 28031 16167
rect 28641 16133 28675 16167
rect 30849 16133 30883 16167
rect 30941 16133 30975 16167
rect 32137 16133 32171 16167
rect 11529 16065 11563 16099
rect 13737 16065 13771 16099
rect 14004 16065 14038 16099
rect 17325 16065 17359 16099
rect 17601 16065 17635 16099
rect 18521 16065 18555 16099
rect 18797 16065 18831 16099
rect 19257 16065 19291 16099
rect 19513 16065 19547 16099
rect 21833 16065 21867 16099
rect 22661 16065 22695 16099
rect 22753 16065 22787 16099
rect 23673 16065 23707 16099
rect 23857 16065 23891 16099
rect 25697 16065 25731 16099
rect 26985 16065 27019 16099
rect 27169 16065 27203 16099
rect 27813 16065 27847 16099
rect 28089 16065 28123 16099
rect 28825 16065 28859 16099
rect 29469 16065 29503 16099
rect 32321 16065 32355 16099
rect 32413 16065 32447 16099
rect 47593 16065 47627 16099
rect 22845 15997 22879 16031
rect 22937 15997 22971 16031
rect 24961 15997 24995 16031
rect 25605 15997 25639 16031
rect 29745 15997 29779 16031
rect 31033 15997 31067 16031
rect 18521 15929 18555 15963
rect 20637 15929 20671 15963
rect 27813 15929 27847 15963
rect 30021 15929 30055 15963
rect 15117 15861 15151 15895
rect 17141 15861 17175 15895
rect 22477 15861 22511 15895
rect 25605 15861 25639 15895
rect 25881 15861 25915 15895
rect 27077 15861 27111 15895
rect 29837 15861 29871 15895
rect 32137 15861 32171 15895
rect 32597 15861 32631 15895
rect 47685 15861 47719 15895
rect 18153 15657 18187 15691
rect 22477 15657 22511 15691
rect 22937 15657 22971 15691
rect 24685 15657 24719 15691
rect 25513 15657 25547 15691
rect 26341 15657 26375 15691
rect 28641 15657 28675 15691
rect 30113 15657 30147 15691
rect 30849 15657 30883 15691
rect 19625 15589 19659 15623
rect 25697 15589 25731 15623
rect 28089 15589 28123 15623
rect 10609 15521 10643 15555
rect 12357 15521 12391 15555
rect 21097 15521 21131 15555
rect 25329 15521 25363 15555
rect 32045 15521 32079 15555
rect 32137 15521 32171 15555
rect 46305 15521 46339 15555
rect 46489 15521 46523 15555
rect 48145 15521 48179 15555
rect 12909 15453 12943 15487
rect 16773 15453 16807 15487
rect 19441 15453 19475 15487
rect 23121 15453 23155 15487
rect 23305 15453 23339 15487
rect 23397 15453 23431 15487
rect 24501 15453 24535 15487
rect 25237 15453 25271 15487
rect 25513 15453 25547 15487
rect 27077 15453 27111 15487
rect 28549 15453 28583 15487
rect 28733 15453 28767 15487
rect 29837 15453 29871 15487
rect 30205 15453 30239 15487
rect 30849 15453 30883 15487
rect 30941 15453 30975 15487
rect 31769 15453 31803 15487
rect 31953 15453 31987 15487
rect 32321 15453 32355 15487
rect 10793 15385 10827 15419
rect 17040 15385 17074 15419
rect 21364 15385 21398 15419
rect 26157 15385 26191 15419
rect 26357 15385 26391 15419
rect 27905 15385 27939 15419
rect 13093 15317 13127 15351
rect 26525 15317 26559 15351
rect 27169 15317 27203 15351
rect 30389 15317 30423 15351
rect 31217 15317 31251 15351
rect 32505 15317 32539 15351
rect 10793 15113 10827 15147
rect 22109 15113 22143 15147
rect 25697 15113 25731 15147
rect 26249 15113 26283 15147
rect 28365 15113 28399 15147
rect 29837 15113 29871 15147
rect 30757 15113 30791 15147
rect 31585 15113 31619 15147
rect 33977 15113 34011 15147
rect 46857 15113 46891 15147
rect 23397 15045 23431 15079
rect 24133 15045 24167 15079
rect 27230 15045 27264 15079
rect 29377 15045 29411 15079
rect 32842 15045 32876 15079
rect 10701 14977 10735 15011
rect 19533 14977 19567 15011
rect 22293 14977 22327 15011
rect 22569 14977 22603 15011
rect 24041 14977 24075 15011
rect 24225 14977 24259 15011
rect 24777 14977 24811 15011
rect 25697 14977 25731 15011
rect 26433 14977 26467 15011
rect 29653 14977 29687 15011
rect 30481 14977 30515 15011
rect 30573 14977 30607 15011
rect 31217 14977 31251 15011
rect 31401 14977 31435 15011
rect 47041 14977 47075 15011
rect 19717 14909 19751 14943
rect 26985 14909 27019 14943
rect 29561 14909 29595 14943
rect 32597 14909 32631 14943
rect 22477 14841 22511 14875
rect 23489 14773 23523 14807
rect 24961 14773 24995 14807
rect 29653 14773 29687 14807
rect 47777 14773 47811 14807
rect 19441 14569 19475 14603
rect 25237 14569 25271 14603
rect 30205 14569 30239 14603
rect 31217 14569 31251 14603
rect 21281 14501 21315 14535
rect 28917 14501 28951 14535
rect 32873 14501 32907 14535
rect 30757 14433 30791 14467
rect 31953 14433 31987 14467
rect 33333 14433 33367 14467
rect 33425 14433 33459 14467
rect 46305 14433 46339 14467
rect 2053 14365 2087 14399
rect 19349 14365 19383 14399
rect 21097 14365 21131 14399
rect 22845 14365 22879 14399
rect 23029 14365 23063 14399
rect 26617 14365 26651 14399
rect 26801 14365 26835 14399
rect 27629 14365 27663 14399
rect 28733 14365 28767 14399
rect 29837 14365 29871 14399
rect 30849 14365 30883 14399
rect 31677 14365 31711 14399
rect 31861 14365 31895 14399
rect 32045 14365 32079 14399
rect 32229 14365 32263 14399
rect 20269 14297 20303 14331
rect 25145 14297 25179 14331
rect 27813 14297 27847 14331
rect 30021 14297 30055 14331
rect 33241 14297 33275 14331
rect 46489 14297 46523 14331
rect 48145 14297 48179 14331
rect 20545 14229 20579 14263
rect 32413 14229 32447 14263
rect 24777 14025 24811 14059
rect 27169 14025 27203 14059
rect 27997 14025 28031 14059
rect 31401 14025 31435 14059
rect 33793 14025 33827 14059
rect 46857 14025 46891 14059
rect 48053 14025 48087 14059
rect 20821 13957 20855 13991
rect 24409 13957 24443 13991
rect 24609 13957 24643 13991
rect 25513 13957 25547 13991
rect 26249 13957 26283 13991
rect 26433 13957 26467 13991
rect 32680 13957 32714 13991
rect 1777 13889 1811 13923
rect 17141 13889 17175 13923
rect 19625 13889 19659 13923
rect 19717 13889 19751 13923
rect 19901 13889 19935 13923
rect 19993 13889 20027 13923
rect 20637 13889 20671 13923
rect 23489 13889 23523 13923
rect 23581 13889 23615 13923
rect 25237 13889 25271 13923
rect 26985 13889 27019 13923
rect 27813 13889 27847 13923
rect 29469 13889 29503 13923
rect 29653 13889 29687 13923
rect 31033 13889 31067 13923
rect 32413 13889 32447 13923
rect 46765 13889 46799 13923
rect 47869 13889 47903 13923
rect 1961 13821 1995 13855
rect 2789 13821 2823 13855
rect 17325 13821 17359 13855
rect 18061 13821 18095 13855
rect 20453 13821 20487 13855
rect 23857 13821 23891 13855
rect 23949 13821 23983 13855
rect 25513 13821 25547 13855
rect 29561 13821 29595 13855
rect 30113 13821 30147 13855
rect 31125 13821 31159 13855
rect 30389 13753 30423 13787
rect 19441 13685 19475 13719
rect 23305 13685 23339 13719
rect 24593 13685 24627 13719
rect 25329 13685 25363 13719
rect 30573 13685 30607 13719
rect 31033 13685 31067 13719
rect 2145 13481 2179 13515
rect 17325 13481 17359 13515
rect 29929 13481 29963 13515
rect 30481 13481 30515 13515
rect 26249 13413 26283 13447
rect 30849 13413 30883 13447
rect 19257 13345 19291 13379
rect 24777 13345 24811 13379
rect 25513 13345 25547 13379
rect 30941 13345 30975 13379
rect 32137 13345 32171 13379
rect 32321 13345 32355 13379
rect 2053 13277 2087 13311
rect 17233 13277 17267 13311
rect 19524 13277 19558 13311
rect 22201 13277 22235 13311
rect 22468 13277 22502 13311
rect 24409 13277 24443 13311
rect 25237 13277 25271 13311
rect 25329 13277 25363 13311
rect 26065 13277 26099 13311
rect 27905 13277 27939 13311
rect 29745 13277 29779 13311
rect 30021 13277 30055 13311
rect 30665 13277 30699 13311
rect 32045 13277 32079 13311
rect 24593 13209 24627 13243
rect 20637 13141 20671 13175
rect 23581 13141 23615 13175
rect 25513 13141 25547 13175
rect 27997 13141 28031 13175
rect 29561 13141 29595 13175
rect 31677 13141 31711 13175
rect 25237 12937 25271 12971
rect 27169 12937 27203 12971
rect 24869 12869 24903 12903
rect 26157 12869 26191 12903
rect 26985 12869 27019 12903
rect 29009 12869 29043 12903
rect 29929 12869 29963 12903
rect 36645 12869 36679 12903
rect 37473 12869 37507 12903
rect 1685 12801 1719 12835
rect 16865 12801 16899 12835
rect 18245 12801 18279 12835
rect 18521 12801 18555 12835
rect 20821 12801 20855 12835
rect 21005 12801 21039 12835
rect 22017 12801 22051 12835
rect 22201 12801 22235 12835
rect 22845 12801 22879 12835
rect 22937 12801 22971 12835
rect 23213 12801 23247 12835
rect 24041 12801 24075 12835
rect 25053 12801 25087 12835
rect 25329 12801 25363 12835
rect 25789 12801 25823 12835
rect 25937 12801 25971 12835
rect 26065 12801 26099 12835
rect 26254 12801 26288 12835
rect 27261 12801 27295 12835
rect 29653 12801 29687 12835
rect 29837 12801 29871 12835
rect 30021 12801 30055 12835
rect 36553 12801 36587 12835
rect 1409 12733 1443 12767
rect 19533 12733 19567 12767
rect 19809 12733 19843 12767
rect 22109 12733 22143 12767
rect 23121 12733 23155 12767
rect 24133 12733 24167 12767
rect 24317 12733 24351 12767
rect 37289 12733 37323 12767
rect 39129 12733 39163 12767
rect 26985 12665 27019 12699
rect 16957 12597 16991 12631
rect 21189 12597 21223 12631
rect 22661 12597 22695 12631
rect 23673 12597 23707 12631
rect 26433 12597 26467 12631
rect 29101 12597 29135 12631
rect 30205 12597 30239 12631
rect 21189 12393 21223 12427
rect 24685 12393 24719 12427
rect 25145 12393 25179 12427
rect 29561 12393 29595 12427
rect 23765 12325 23799 12359
rect 22937 12257 22971 12291
rect 23121 12257 23155 12291
rect 24869 12257 24903 12291
rect 18521 12189 18555 12223
rect 19809 12189 19843 12223
rect 23673 12189 23707 12223
rect 23857 12189 23891 12223
rect 24961 12189 24995 12223
rect 26157 12189 26191 12223
rect 28273 12189 28307 12223
rect 29745 12189 29779 12223
rect 29837 12189 29871 12223
rect 30021 12189 30055 12223
rect 30113 12189 30147 12223
rect 18705 12121 18739 12155
rect 20076 12121 20110 12155
rect 24685 12121 24719 12155
rect 26424 12121 26458 12155
rect 28089 12121 28123 12155
rect 22477 12053 22511 12087
rect 22845 12053 22879 12087
rect 27537 12053 27571 12087
rect 20177 11849 20211 11883
rect 23949 11849 23983 11883
rect 26065 11849 26099 11883
rect 28457 11849 28491 11883
rect 29469 11849 29503 11883
rect 16957 11781 16991 11815
rect 2237 11713 2271 11747
rect 2881 11713 2915 11747
rect 19349 11713 19383 11747
rect 19438 11713 19472 11747
rect 19533 11713 19567 11747
rect 19717 11713 19751 11747
rect 20407 11713 20441 11747
rect 20545 11713 20579 11747
rect 20637 11713 20671 11747
rect 20821 11713 20855 11747
rect 22109 11713 22143 11747
rect 24317 11713 24351 11747
rect 28273 11713 28307 11747
rect 28549 11713 28583 11747
rect 29009 11713 29043 11747
rect 29285 11713 29319 11747
rect 30573 11713 30607 11747
rect 16773 11645 16807 11679
rect 18153 11645 18187 11679
rect 24409 11645 24443 11679
rect 24593 11645 24627 11679
rect 26157 11645 26191 11679
rect 26341 11645 26375 11679
rect 29101 11645 29135 11679
rect 30665 11645 30699 11679
rect 30757 11645 30791 11679
rect 25697 11577 25731 11611
rect 2329 11509 2363 11543
rect 2973 11509 3007 11543
rect 19073 11509 19107 11543
rect 21925 11509 21959 11543
rect 28273 11509 28307 11543
rect 29009 11509 29043 11543
rect 30205 11509 30239 11543
rect 47777 11509 47811 11543
rect 18705 11305 18739 11339
rect 19625 11305 19659 11339
rect 22753 11305 22787 11339
rect 24869 11305 24903 11339
rect 25881 11305 25915 11339
rect 27813 11305 27847 11339
rect 28825 11305 28859 11339
rect 32137 11305 32171 11339
rect 25053 11237 25087 11271
rect 1593 11169 1627 11203
rect 3065 11169 3099 11203
rect 24685 11169 24719 11203
rect 30113 11169 30147 11203
rect 30757 11169 30791 11203
rect 46305 11169 46339 11203
rect 1409 11101 1443 11135
rect 17325 11101 17359 11135
rect 17592 11101 17626 11135
rect 19257 11101 19291 11135
rect 19441 11101 19475 11135
rect 21373 11101 21407 11135
rect 21640 11101 21674 11135
rect 24869 11101 24903 11135
rect 25513 11101 25547 11135
rect 27629 11101 27663 11135
rect 27813 11101 27847 11135
rect 28641 11101 28675 11135
rect 28917 11101 28951 11135
rect 29929 11101 29963 11135
rect 31013 11101 31047 11135
rect 24409 11033 24443 11067
rect 25697 11033 25731 11067
rect 46489 11033 46523 11067
rect 48145 11033 48179 11067
rect 27997 10965 28031 10999
rect 28457 10965 28491 10999
rect 29561 10965 29595 10999
rect 30021 10965 30055 10999
rect 29285 10761 29319 10795
rect 31125 10761 31159 10795
rect 46949 10761 46983 10795
rect 27169 10693 27203 10727
rect 1409 10625 1443 10659
rect 1685 10625 1719 10659
rect 19303 10625 19337 10659
rect 19438 10628 19472 10662
rect 19533 10625 19567 10659
rect 19717 10625 19751 10659
rect 24041 10625 24075 10659
rect 26157 10625 26191 10659
rect 26249 10625 26283 10659
rect 26985 10625 27019 10659
rect 27261 10625 27295 10659
rect 28825 10625 28859 10659
rect 29094 10625 29128 10659
rect 29745 10625 29779 10659
rect 29929 10625 29963 10659
rect 30297 10625 30331 10659
rect 31033 10625 31067 10659
rect 46857 10625 46891 10659
rect 47777 10625 47811 10659
rect 2881 10557 2915 10591
rect 24501 10557 24535 10591
rect 26433 10557 26467 10591
rect 29009 10557 29043 10591
rect 30021 10557 30055 10591
rect 30113 10557 30147 10591
rect 26985 10489 27019 10523
rect 47961 10489 47995 10523
rect 3525 10421 3559 10455
rect 19073 10421 19107 10455
rect 24317 10421 24351 10455
rect 26341 10421 26375 10455
rect 28825 10421 28859 10455
rect 30481 10421 30515 10455
rect 19625 10217 19659 10251
rect 24409 10217 24443 10251
rect 26065 10217 26099 10251
rect 28457 10217 28491 10251
rect 29929 10217 29963 10251
rect 31953 10217 31987 10251
rect 1409 10081 1443 10115
rect 23406 10081 23440 10115
rect 24869 10081 24903 10115
rect 25053 10081 25087 10115
rect 26525 10081 26559 10115
rect 26709 10081 26743 10115
rect 28641 10081 28675 10115
rect 19257 10013 19291 10047
rect 20545 10013 20579 10047
rect 20637 10013 20671 10047
rect 20729 10013 20763 10047
rect 20913 10013 20947 10047
rect 23121 10013 23155 10047
rect 23305 10013 23339 10047
rect 23489 10013 23523 10047
rect 23673 10013 23707 10047
rect 24777 10013 24811 10047
rect 28365 10013 28399 10047
rect 29561 10013 29595 10047
rect 30573 10013 30607 10047
rect 30840 10013 30874 10047
rect 1593 9945 1627 9979
rect 3249 9945 3283 9979
rect 19441 9945 19475 9979
rect 29745 9945 29779 9979
rect 20269 9877 20303 9911
rect 23857 9877 23891 9911
rect 26433 9877 26467 9911
rect 28917 9877 28951 9911
rect 20821 9673 20855 9707
rect 24501 9673 24535 9707
rect 29653 9673 29687 9707
rect 17877 9537 17911 9571
rect 18144 9537 18178 9571
rect 20453 9537 20487 9571
rect 20637 9537 20671 9571
rect 23121 9537 23155 9571
rect 23388 9537 23422 9571
rect 25697 9537 25731 9571
rect 25881 9537 25915 9571
rect 26249 9537 26283 9571
rect 28365 9537 28399 9571
rect 29469 9537 29503 9571
rect 29653 9537 29687 9571
rect 25973 9469 26007 9503
rect 26065 9469 26099 9503
rect 28457 9469 28491 9503
rect 28549 9469 28583 9503
rect 27997 9401 28031 9435
rect 19257 9333 19291 9367
rect 26433 9333 26467 9367
rect 27353 9129 27387 9163
rect 17325 8993 17359 9027
rect 25973 8993 26007 9027
rect 28457 8993 28491 9027
rect 19809 8925 19843 8959
rect 19901 8925 19935 8959
rect 19993 8925 20027 8959
rect 20177 8925 20211 8959
rect 20637 8925 20671 8959
rect 20904 8925 20938 8959
rect 26240 8925 26274 8959
rect 28181 8925 28215 8959
rect 28365 8925 28399 8959
rect 28549 8925 28583 8959
rect 28733 8925 28767 8959
rect 17592 8857 17626 8891
rect 19533 8857 19567 8891
rect 47961 8857 47995 8891
rect 18705 8789 18739 8823
rect 22017 8789 22051 8823
rect 28917 8789 28951 8823
rect 48053 8789 48087 8823
rect 29745 8585 29779 8619
rect 47869 8585 47903 8619
rect 1869 8449 1903 8483
rect 18521 8449 18555 8483
rect 28365 8449 28399 8483
rect 28632 8449 28666 8483
rect 30481 8449 30515 8483
rect 30573 8449 30607 8483
rect 30665 8449 30699 8483
rect 30849 8449 30883 8483
rect 47777 8449 47811 8483
rect 18705 8381 18739 8415
rect 19441 8381 19475 8415
rect 2145 8313 2179 8347
rect 30205 8245 30239 8279
rect 18613 8041 18647 8075
rect 19809 8041 19843 8075
rect 31861 8041 31895 8075
rect 24777 7905 24811 7939
rect 28089 7905 28123 7939
rect 18521 7837 18555 7871
rect 19625 7837 19659 7871
rect 21189 7837 21223 7871
rect 21278 7837 21312 7871
rect 21373 7837 21407 7871
rect 21557 7837 21591 7871
rect 22017 7837 22051 7871
rect 22201 7837 22235 7871
rect 23489 7837 23523 7871
rect 23581 7837 23615 7871
rect 23673 7837 23707 7871
rect 23857 7837 23891 7871
rect 24593 7837 24627 7871
rect 26893 7837 26927 7871
rect 26985 7837 27019 7871
rect 27077 7837 27111 7871
rect 27261 7837 27295 7871
rect 29653 7837 29687 7871
rect 31493 7837 31527 7871
rect 1869 7769 1903 7803
rect 19441 7769 19475 7803
rect 24409 7769 24443 7803
rect 27721 7769 27755 7803
rect 27905 7769 27939 7803
rect 29920 7769 29954 7803
rect 31677 7769 31711 7803
rect 2145 7701 2179 7735
rect 20913 7701 20947 7735
rect 22385 7701 22419 7735
rect 23213 7701 23247 7735
rect 26617 7701 26651 7735
rect 31033 7701 31067 7735
rect 23213 7497 23247 7531
rect 27230 7429 27264 7463
rect 18889 7361 18923 7395
rect 22089 7361 22123 7395
rect 23929 7361 23963 7395
rect 26249 7361 26283 7395
rect 29653 7361 29687 7395
rect 46673 7361 46707 7395
rect 19073 7293 19107 7327
rect 19441 7293 19475 7327
rect 21833 7293 21867 7327
rect 23673 7293 23707 7327
rect 26985 7293 27019 7327
rect 29837 7293 29871 7327
rect 30113 7293 30147 7327
rect 2053 7157 2087 7191
rect 25053 7157 25087 7191
rect 26341 7157 26375 7191
rect 28365 7157 28399 7191
rect 46765 7157 46799 7191
rect 47777 7157 47811 7191
rect 22477 6953 22511 6987
rect 25789 6953 25823 6987
rect 29837 6953 29871 6987
rect 1409 6817 1443 6851
rect 2789 6817 2823 6851
rect 19349 6817 19383 6851
rect 19993 6817 20027 6851
rect 21097 6817 21131 6851
rect 23213 6817 23247 6851
rect 26709 6817 26743 6851
rect 26985 6817 27019 6851
rect 46489 6817 46523 6851
rect 48145 6817 48179 6851
rect 19257 6749 19291 6783
rect 20269 6749 20303 6783
rect 20361 6749 20395 6783
rect 20453 6749 20487 6783
rect 20637 6749 20671 6783
rect 21353 6749 21387 6783
rect 23443 6749 23477 6783
rect 23581 6749 23615 6783
rect 23673 6749 23707 6783
rect 23857 6749 23891 6783
rect 24409 6749 24443 6783
rect 26525 6749 26559 6783
rect 29745 6749 29779 6783
rect 46305 6749 46339 6783
rect 1593 6681 1627 6715
rect 24654 6681 24688 6715
rect 2237 6409 2271 6443
rect 22201 6409 22235 6443
rect 23489 6409 23523 6443
rect 22017 6341 22051 6375
rect 23305 6341 23339 6375
rect 2145 6273 2179 6307
rect 21833 6273 21867 6307
rect 23121 6273 23155 6307
rect 24685 5865 24719 5899
rect 25053 5865 25087 5899
rect 25513 5865 25547 5899
rect 25237 5729 25271 5763
rect 48145 5729 48179 5763
rect 2329 5661 2363 5695
rect 2973 5661 3007 5695
rect 25329 5661 25363 5695
rect 47409 5661 47443 5695
rect 25053 5593 25087 5627
rect 47961 5593 47995 5627
rect 3065 5525 3099 5559
rect 2329 5253 2363 5287
rect 2145 5185 2179 5219
rect 46857 5185 46891 5219
rect 47593 5185 47627 5219
rect 2789 5117 2823 5151
rect 1685 4981 1719 5015
rect 46949 4981 46983 5015
rect 47685 4981 47719 5015
rect 1409 4641 1443 4675
rect 1593 4641 1627 4675
rect 3893 4641 3927 4675
rect 22017 4641 22051 4675
rect 41889 4641 41923 4675
rect 43269 4641 43303 4675
rect 46305 4641 46339 4675
rect 46489 4641 46523 4675
rect 48145 4641 48179 4675
rect 3249 4573 3283 4607
rect 3801 4573 3835 4607
rect 6285 4573 6319 4607
rect 6929 4573 6963 4607
rect 8033 4573 8067 4607
rect 30481 4573 30515 4607
rect 31125 4573 31159 4607
rect 45201 4573 45235 4607
rect 45845 4573 45879 4607
rect 22201 4505 22235 4539
rect 23857 4505 23891 4539
rect 42073 4505 42107 4539
rect 8125 4437 8159 4471
rect 22661 4233 22695 4267
rect 42533 4233 42567 4267
rect 8125 4165 8159 4199
rect 47961 4165 47995 4199
rect 2053 4097 2087 4131
rect 2697 4097 2731 4131
rect 6377 4097 6411 4131
rect 7021 4097 7055 4131
rect 7941 4097 7975 4131
rect 11621 4097 11655 4131
rect 12541 4097 12575 4131
rect 22569 4097 22603 4131
rect 30757 4097 30791 4131
rect 31401 4097 31435 4131
rect 36369 4097 36403 4131
rect 37841 4097 37875 4131
rect 40969 4097 41003 4131
rect 42441 4097 42475 4131
rect 43453 4097 43487 4131
rect 46397 4097 46431 4131
rect 8401 4029 8435 4063
rect 13185 4029 13219 4063
rect 13369 4029 13403 4063
rect 13645 4029 13679 4063
rect 44097 4029 44131 4063
rect 44281 4029 44315 4063
rect 44557 4029 44591 4063
rect 12633 3961 12667 3995
rect 43545 3961 43579 3995
rect 1593 3893 1627 3927
rect 2145 3893 2179 3927
rect 2789 3893 2823 3927
rect 3801 3893 3835 3927
rect 5457 3893 5491 3927
rect 6469 3893 6503 3927
rect 7113 3893 7147 3927
rect 11713 3893 11747 3927
rect 17601 3893 17635 3927
rect 21005 3893 21039 3927
rect 23673 3893 23707 3927
rect 25973 3893 26007 3927
rect 30021 3893 30055 3927
rect 30849 3893 30883 3927
rect 31493 3893 31527 3927
rect 32413 3893 32447 3927
rect 36461 3893 36495 3927
rect 37933 3893 37967 3927
rect 41061 3893 41095 3927
rect 41797 3893 41831 3927
rect 46489 3893 46523 3927
rect 48053 3893 48087 3927
rect 22661 3689 22695 3723
rect 43085 3689 43119 3723
rect 43821 3689 43855 3723
rect 1593 3553 1627 3587
rect 1869 3553 1903 3587
rect 5181 3553 5215 3587
rect 5365 3553 5399 3587
rect 6561 3553 6595 3587
rect 12817 3553 12851 3587
rect 20729 3553 20763 3587
rect 25697 3553 25731 3587
rect 26433 3553 26467 3587
rect 30849 3553 30883 3587
rect 31033 3553 31067 3587
rect 31585 3553 31619 3587
rect 36277 3553 36311 3587
rect 36737 3553 36771 3587
rect 40785 3553 40819 3587
rect 41245 3553 41279 3587
rect 44465 3553 44499 3587
rect 46029 3553 46063 3587
rect 46213 3553 46247 3587
rect 46489 3553 46523 3587
rect 1409 3485 1443 3519
rect 4353 3485 4387 3519
rect 7481 3485 7515 3519
rect 11713 3485 11747 3519
rect 14473 3485 14507 3519
rect 15117 3485 15151 3519
rect 17693 3485 17727 3519
rect 19625 3485 19659 3519
rect 20269 3485 20303 3519
rect 22845 3485 22879 3519
rect 23305 3485 23339 3519
rect 29561 3485 29595 3519
rect 30205 3485 30239 3519
rect 36093 3485 36127 3519
rect 38761 3485 38795 3519
rect 39957 3485 39991 3519
rect 40601 3485 40635 3519
rect 45017 3485 45051 3519
rect 7573 3417 7607 3451
rect 11897 3417 11931 3451
rect 14565 3417 14599 3451
rect 15301 3417 15335 3451
rect 16957 3417 16991 3451
rect 19717 3417 19751 3451
rect 20453 3417 20487 3451
rect 25881 3417 25915 3451
rect 4445 3349 4479 3383
rect 17785 3349 17819 3383
rect 23397 3349 23431 3383
rect 29653 3349 29687 3383
rect 30297 3349 30331 3383
rect 45109 3349 45143 3383
rect 1961 3145 1995 3179
rect 1869 3077 1903 3111
rect 3709 3077 3743 3111
rect 17509 3077 17543 3111
rect 23581 3077 23615 3111
rect 29926 3077 29960 3111
rect 32321 3077 32355 3111
rect 44925 3077 44959 3111
rect 2605 3009 2639 3043
rect 3525 3009 3559 3043
rect 6377 3009 6411 3043
rect 10057 3009 10091 3043
rect 10241 3009 10275 3043
rect 11989 3009 12023 3043
rect 15301 3009 15335 3043
rect 17325 3009 17359 3043
rect 20453 3009 20487 3043
rect 22753 3009 22787 3043
rect 23397 3009 23431 3043
rect 26065 3009 26099 3043
rect 29745 3009 29779 3043
rect 32137 3009 32171 3043
rect 36277 3009 36311 3043
rect 38577 3009 38611 3043
rect 41521 3009 41555 3043
rect 42441 3009 42475 3043
rect 44741 3009 44775 3043
rect 47869 3009 47903 3043
rect 2789 2941 2823 2975
rect 3985 2941 4019 2975
rect 6561 2941 6595 2975
rect 6837 2941 6871 2975
rect 8677 2941 8711 2975
rect 8953 2941 8987 2975
rect 12449 2941 12483 2975
rect 12633 2941 12667 2975
rect 12909 2941 12943 2975
rect 18061 2941 18095 2975
rect 23857 2941 23891 2975
rect 31309 2941 31343 2975
rect 33517 2941 33551 2975
rect 38761 2941 38795 2975
rect 39957 2941 39991 2975
rect 41613 2941 41647 2975
rect 42625 2941 42659 2975
rect 42901 2941 42935 2975
rect 45201 2941 45235 2975
rect 48053 2873 48087 2907
rect 22845 2805 22879 2839
rect 26157 2805 26191 2839
rect 3985 2601 4019 2635
rect 12725 2601 12759 2635
rect 13369 2601 13403 2635
rect 17785 2533 17819 2567
rect 20361 2533 20395 2567
rect 25881 2533 25915 2567
rect 27261 2533 27295 2567
rect 33149 2533 33183 2567
rect 35081 2533 35115 2567
rect 36185 2533 36219 2567
rect 1409 2465 1443 2499
rect 1869 2465 1903 2499
rect 6377 2465 6411 2499
rect 6561 2465 6595 2499
rect 7021 2465 7055 2499
rect 8953 2465 8987 2499
rect 9229 2465 9263 2499
rect 21833 2465 21867 2499
rect 22293 2465 22327 2499
rect 24869 2465 24903 2499
rect 28089 2465 28123 2499
rect 29745 2465 29779 2499
rect 29929 2465 29963 2499
rect 30941 2465 30975 2499
rect 38761 2465 38795 2499
rect 45201 2465 45235 2499
rect 4629 2397 4663 2431
rect 14749 2397 14783 2431
rect 24593 2397 24627 2431
rect 26065 2397 26099 2431
rect 27077 2397 27111 2431
rect 27813 2397 27847 2431
rect 32965 2397 32999 2431
rect 34897 2397 34931 2431
rect 36369 2397 36403 2431
rect 38485 2397 38519 2431
rect 44465 2397 44499 2431
rect 47041 2397 47075 2431
rect 1593 2329 1627 2363
rect 10333 2329 10367 2363
rect 14565 2329 14599 2363
rect 17601 2329 17635 2363
rect 20177 2329 20211 2363
rect 22017 2329 22051 2363
rect 33977 2329 34011 2363
rect 43361 2329 43395 2363
rect 44281 2329 44315 2363
rect 45385 2329 45419 2363
rect 47777 2329 47811 2363
rect 4813 2261 4847 2295
rect 10609 2261 10643 2295
rect 34069 2261 34103 2295
rect 43453 2261 43487 2295
rect 47869 2261 47903 2295
<< metal1 >>
rect 4062 49716 4068 49768
rect 4120 49756 4126 49768
rect 5626 49756 5632 49768
rect 4120 49728 5632 49756
rect 4120 49716 4126 49728
rect 5626 49716 5632 49728
rect 5684 49716 5690 49768
rect 36998 49716 37004 49768
rect 37056 49756 37062 49768
rect 45554 49756 45560 49768
rect 37056 49728 45560 49756
rect 37056 49716 37062 49728
rect 45554 49716 45560 49728
rect 45612 49716 45618 49768
rect 1104 49530 48852 49552
rect 1104 49478 4214 49530
rect 4266 49478 4278 49530
rect 4330 49478 4342 49530
rect 4394 49478 4406 49530
rect 4458 49478 4470 49530
rect 4522 49478 34934 49530
rect 34986 49478 34998 49530
rect 35050 49478 35062 49530
rect 35114 49478 35126 49530
rect 35178 49478 35190 49530
rect 35242 49478 48852 49530
rect 1104 49456 48852 49478
rect 24118 49348 24124 49360
rect 22066 49320 24124 49348
rect 6549 49283 6607 49289
rect 6549 49249 6561 49283
rect 6595 49280 6607 49283
rect 6914 49280 6920 49292
rect 6595 49252 6920 49280
rect 6595 49249 6607 49252
rect 6549 49243 6607 49249
rect 6914 49240 6920 49252
rect 6972 49240 6978 49292
rect 7098 49280 7104 49292
rect 7059 49252 7104 49280
rect 7098 49240 7104 49252
rect 7156 49240 7162 49292
rect 7742 49240 7748 49292
rect 7800 49280 7806 49292
rect 9401 49283 9459 49289
rect 9401 49280 9413 49283
rect 7800 49252 9413 49280
rect 7800 49240 7806 49252
rect 9401 49249 9413 49252
rect 9447 49249 9459 49283
rect 12710 49280 12716 49292
rect 12671 49252 12716 49280
rect 9401 49243 9459 49249
rect 12710 49240 12716 49252
rect 12768 49240 12774 49292
rect 14458 49240 14464 49292
rect 14516 49280 14522 49292
rect 14516 49252 15424 49280
rect 14516 49240 14522 49252
rect 658 49172 664 49224
rect 716 49212 722 49224
rect 1857 49215 1915 49221
rect 1857 49212 1869 49215
rect 716 49184 1869 49212
rect 716 49172 722 49184
rect 1857 49181 1869 49184
rect 1903 49181 1915 49215
rect 1857 49175 1915 49181
rect 3602 49172 3608 49224
rect 3660 49212 3666 49224
rect 4249 49215 4307 49221
rect 4249 49212 4261 49215
rect 3660 49184 4261 49212
rect 3660 49172 3666 49184
rect 4249 49181 4261 49184
rect 4295 49181 4307 49215
rect 4249 49175 4307 49181
rect 4614 49172 4620 49224
rect 4672 49212 4678 49224
rect 5077 49215 5135 49221
rect 5077 49212 5089 49215
rect 4672 49184 5089 49212
rect 4672 49172 4678 49184
rect 5077 49181 5089 49184
rect 5123 49181 5135 49215
rect 8938 49212 8944 49224
rect 8899 49184 8944 49212
rect 5077 49175 5135 49181
rect 8938 49172 8944 49184
rect 8996 49172 9002 49224
rect 11606 49172 11612 49224
rect 11664 49212 11670 49224
rect 11977 49215 12035 49221
rect 11977 49212 11989 49215
rect 11664 49184 11989 49212
rect 11664 49172 11670 49184
rect 11977 49181 11989 49184
rect 12023 49181 12035 49215
rect 11977 49175 12035 49181
rect 12989 49215 13047 49221
rect 12989 49181 13001 49215
rect 13035 49181 13047 49215
rect 12989 49175 13047 49181
rect 2774 49144 2780 49156
rect 2735 49116 2780 49144
rect 2774 49104 2780 49116
rect 2832 49104 2838 49156
rect 2958 49144 2964 49156
rect 2919 49116 2964 49144
rect 2958 49104 2964 49116
rect 3016 49104 3022 49156
rect 6733 49147 6791 49153
rect 6733 49113 6745 49147
rect 6779 49144 6791 49147
rect 7374 49144 7380 49156
rect 6779 49116 7380 49144
rect 6779 49113 6791 49116
rect 6733 49107 6791 49113
rect 7374 49104 7380 49116
rect 7432 49104 7438 49156
rect 8478 49104 8484 49156
rect 8536 49144 8542 49156
rect 9125 49147 9183 49153
rect 9125 49144 9137 49147
rect 8536 49116 9137 49144
rect 8536 49104 8542 49116
rect 9125 49113 9137 49116
rect 9171 49113 9183 49147
rect 13004 49144 13032 49175
rect 13814 49172 13820 49224
rect 13872 49212 13878 49224
rect 15396 49221 15424 49252
rect 16574 49240 16580 49292
rect 16632 49280 16638 49292
rect 16669 49283 16727 49289
rect 16669 49280 16681 49283
rect 16632 49252 16681 49280
rect 16632 49240 16638 49252
rect 16669 49249 16681 49252
rect 16715 49249 16727 49283
rect 16669 49243 16727 49249
rect 16945 49283 17003 49289
rect 16945 49249 16957 49283
rect 16991 49280 17003 49283
rect 22066 49280 22094 49320
rect 24118 49308 24124 49320
rect 24176 49308 24182 49360
rect 28997 49351 29055 49357
rect 28997 49317 29009 49351
rect 29043 49348 29055 49351
rect 29914 49348 29920 49360
rect 29043 49320 29920 49348
rect 29043 49317 29055 49320
rect 28997 49311 29055 49317
rect 29914 49308 29920 49320
rect 29972 49308 29978 49360
rect 33502 49308 33508 49360
rect 33560 49348 33566 49360
rect 34422 49348 34428 49360
rect 33560 49320 34428 49348
rect 33560 49308 33566 49320
rect 34422 49308 34428 49320
rect 34480 49308 34486 49360
rect 22554 49280 22560 49292
rect 16991 49252 22094 49280
rect 22515 49252 22560 49280
rect 16991 49249 17003 49252
rect 16945 49243 17003 49249
rect 22554 49240 22560 49252
rect 22612 49240 22618 49292
rect 29733 49283 29791 49289
rect 29733 49249 29745 49283
rect 29779 49280 29791 49283
rect 30466 49280 30472 49292
rect 29779 49252 30472 49280
rect 29779 49249 29791 49252
rect 29733 49243 29791 49249
rect 30466 49240 30472 49252
rect 30524 49240 30530 49292
rect 30926 49280 30932 49292
rect 30887 49252 30932 49280
rect 30926 49240 30932 49252
rect 30984 49240 30990 49292
rect 43162 49280 43168 49292
rect 43123 49252 43168 49280
rect 43162 49240 43168 49252
rect 43220 49240 43226 49292
rect 45186 49240 45192 49292
rect 45244 49280 45250 49292
rect 45557 49283 45615 49289
rect 45557 49280 45569 49283
rect 45244 49252 45569 49280
rect 45244 49240 45250 49252
rect 45557 49249 45569 49252
rect 45603 49249 45615 49283
rect 45557 49243 45615 49249
rect 14553 49215 14611 49221
rect 14553 49212 14565 49215
rect 13872 49184 14565 49212
rect 13872 49172 13878 49184
rect 14553 49181 14565 49184
rect 14599 49181 14611 49215
rect 14553 49175 14611 49181
rect 15381 49215 15439 49221
rect 15381 49181 15393 49215
rect 15427 49181 15439 49215
rect 15381 49175 15439 49181
rect 17954 49172 17960 49224
rect 18012 49212 18018 49224
rect 18141 49215 18199 49221
rect 18141 49212 18153 49215
rect 18012 49184 18153 49212
rect 18012 49172 18018 49184
rect 18141 49181 18153 49184
rect 18187 49181 18199 49215
rect 19426 49212 19432 49224
rect 19387 49184 19432 49212
rect 18141 49175 18199 49181
rect 19426 49172 19432 49184
rect 19484 49172 19490 49224
rect 20070 49212 20076 49224
rect 20031 49184 20076 49212
rect 20070 49172 20076 49184
rect 20128 49172 20134 49224
rect 21269 49215 21327 49221
rect 21269 49181 21281 49215
rect 21315 49212 21327 49215
rect 21634 49212 21640 49224
rect 21315 49184 21640 49212
rect 21315 49181 21327 49184
rect 21269 49175 21327 49181
rect 21634 49172 21640 49184
rect 21692 49172 21698 49224
rect 21818 49212 21824 49224
rect 21779 49184 21824 49212
rect 21818 49172 21824 49184
rect 21876 49172 21882 49224
rect 23842 49172 23848 49224
rect 23900 49212 23906 49224
rect 24581 49215 24639 49221
rect 24581 49212 24593 49215
rect 23900 49184 24593 49212
rect 23900 49172 23906 49184
rect 24581 49181 24593 49184
rect 24627 49181 24639 49215
rect 25958 49212 25964 49224
rect 25919 49184 25964 49212
rect 24581 49175 24639 49181
rect 25958 49172 25964 49184
rect 26016 49172 26022 49224
rect 26418 49172 26424 49224
rect 26476 49212 26482 49224
rect 27433 49215 27491 49221
rect 27433 49212 27445 49215
rect 26476 49184 27445 49212
rect 26476 49172 26482 49184
rect 27433 49181 27445 49184
rect 27479 49181 27491 49215
rect 27433 49175 27491 49181
rect 27982 49172 27988 49224
rect 28040 49212 28046 49224
rect 28261 49215 28319 49221
rect 28261 49212 28273 49215
rect 28040 49184 28273 49212
rect 28040 49172 28046 49184
rect 28261 49181 28273 49184
rect 28307 49181 28319 49215
rect 28261 49175 28319 49181
rect 28813 49215 28871 49221
rect 28813 49181 28825 49215
rect 28859 49212 28871 49215
rect 28994 49212 29000 49224
rect 28859 49184 29000 49212
rect 28859 49181 28871 49184
rect 28813 49175 28871 49181
rect 28994 49172 29000 49184
rect 29052 49172 29058 49224
rect 31938 49172 31944 49224
rect 31996 49212 32002 49224
rect 33045 49215 33103 49221
rect 33045 49212 33057 49215
rect 31996 49184 33057 49212
rect 31996 49172 32002 49184
rect 33045 49181 33057 49184
rect 33091 49181 33103 49215
rect 33045 49175 33103 49181
rect 33502 49172 33508 49224
rect 33560 49212 33566 49224
rect 33781 49215 33839 49221
rect 33781 49212 33793 49215
rect 33560 49184 33793 49212
rect 33560 49172 33566 49184
rect 33781 49181 33793 49184
rect 33827 49181 33839 49215
rect 33781 49175 33839 49181
rect 34882 49172 34888 49224
rect 34940 49212 34946 49224
rect 35529 49215 35587 49221
rect 35529 49212 35541 49215
rect 34940 49184 35541 49212
rect 34940 49172 34946 49184
rect 35529 49181 35541 49184
rect 35575 49181 35587 49215
rect 36170 49212 36176 49224
rect 36131 49184 36176 49212
rect 35529 49175 35587 49181
rect 36170 49172 36176 49184
rect 36228 49172 36234 49224
rect 38194 49212 38200 49224
rect 38155 49184 38200 49212
rect 38194 49172 38200 49184
rect 38252 49172 38258 49224
rect 40221 49215 40279 49221
rect 40221 49181 40233 49215
rect 40267 49212 40279 49215
rect 42613 49215 42671 49221
rect 42613 49212 42625 49215
rect 40267 49184 42625 49212
rect 40267 49181 40279 49184
rect 40221 49175 40279 49181
rect 42613 49181 42625 49184
rect 42659 49181 42671 49215
rect 42613 49175 42671 49181
rect 43990 49172 43996 49224
rect 44048 49212 44054 49224
rect 45005 49215 45063 49221
rect 45005 49212 45017 49215
rect 44048 49184 45017 49212
rect 44048 49172 44054 49184
rect 45005 49181 45017 49184
rect 45051 49181 45063 49215
rect 47762 49212 47768 49224
rect 47723 49184 47768 49212
rect 45005 49175 45063 49181
rect 47762 49172 47768 49184
rect 47820 49172 47826 49224
rect 17218 49144 17224 49156
rect 13004 49116 17224 49144
rect 9125 49107 9183 49113
rect 17218 49104 17224 49116
rect 17276 49104 17282 49156
rect 19613 49147 19671 49153
rect 19613 49113 19625 49147
rect 19659 49144 19671 49147
rect 20530 49144 20536 49156
rect 19659 49116 20536 49144
rect 19659 49113 19671 49116
rect 19613 49107 19671 49113
rect 20530 49104 20536 49116
rect 20588 49104 20594 49156
rect 22005 49147 22063 49153
rect 22005 49113 22017 49147
rect 22051 49144 22063 49147
rect 22278 49144 22284 49156
rect 22051 49116 22284 49144
rect 22051 49113 22063 49116
rect 22005 49107 22063 49113
rect 22278 49104 22284 49116
rect 22336 49104 22342 49156
rect 27617 49147 27675 49153
rect 27617 49113 27629 49147
rect 27663 49144 27675 49147
rect 27706 49144 27712 49156
rect 27663 49116 27712 49144
rect 27663 49113 27675 49116
rect 27617 49107 27675 49113
rect 27706 49104 27712 49116
rect 27764 49104 27770 49156
rect 29917 49147 29975 49153
rect 29917 49113 29929 49147
rect 29963 49144 29975 49147
rect 30650 49144 30656 49156
rect 29963 49116 30656 49144
rect 29963 49113 29975 49116
rect 29917 49107 29975 49113
rect 30650 49104 30656 49116
rect 30708 49104 30714 49156
rect 40770 49144 40776 49156
rect 40731 49116 40776 49144
rect 40770 49104 40776 49116
rect 40828 49104 40834 49156
rect 41509 49147 41567 49153
rect 41509 49113 41521 49147
rect 41555 49144 41567 49147
rect 41690 49144 41696 49156
rect 41555 49116 41696 49144
rect 41555 49113 41567 49116
rect 41509 49107 41567 49113
rect 41690 49104 41696 49116
rect 41748 49104 41754 49156
rect 41782 49104 41788 49156
rect 41840 49144 41846 49156
rect 42797 49147 42855 49153
rect 42797 49144 42809 49147
rect 41840 49116 42809 49144
rect 41840 49104 41846 49116
rect 42797 49113 42809 49116
rect 42843 49113 42855 49147
rect 42797 49107 42855 49113
rect 44082 49104 44088 49156
rect 44140 49144 44146 49156
rect 45189 49147 45247 49153
rect 45189 49144 45201 49147
rect 44140 49116 45201 49144
rect 44140 49104 44146 49116
rect 45189 49113 45201 49116
rect 45235 49113 45247 49147
rect 45189 49107 45247 49113
rect 1486 49036 1492 49088
rect 1544 49076 1550 49088
rect 1949 49079 2007 49085
rect 1949 49076 1961 49079
rect 1544 49048 1961 49076
rect 1544 49036 1550 49048
rect 1949 49045 1961 49048
rect 1995 49045 2007 49079
rect 1949 49039 2007 49045
rect 4525 49079 4583 49085
rect 4525 49045 4537 49079
rect 4571 49076 4583 49079
rect 4614 49076 4620 49088
rect 4571 49048 4620 49076
rect 4571 49045 4583 49048
rect 4525 49039 4583 49045
rect 4614 49036 4620 49048
rect 4672 49036 4678 49088
rect 5258 49076 5264 49088
rect 5219 49048 5264 49076
rect 5258 49036 5264 49048
rect 5316 49036 5322 49088
rect 12066 49076 12072 49088
rect 12027 49048 12072 49076
rect 12066 49036 12072 49048
rect 12124 49036 12130 49088
rect 14642 49076 14648 49088
rect 14603 49048 14648 49076
rect 14642 49036 14648 49048
rect 14700 49036 14706 49088
rect 15197 49079 15255 49085
rect 15197 49045 15209 49079
rect 15243 49076 15255 49079
rect 17586 49076 17592 49088
rect 15243 49048 17592 49076
rect 15243 49045 15255 49048
rect 15197 49039 15255 49045
rect 17586 49036 17592 49048
rect 17644 49036 17650 49088
rect 20257 49079 20315 49085
rect 20257 49045 20269 49079
rect 20303 49076 20315 49079
rect 20346 49076 20352 49088
rect 20303 49048 20352 49076
rect 20303 49045 20315 49048
rect 20257 49039 20315 49045
rect 20346 49036 20352 49048
rect 20404 49036 20410 49088
rect 21082 49076 21088 49088
rect 21043 49048 21088 49076
rect 21082 49036 21088 49048
rect 21140 49036 21146 49088
rect 22370 49036 22376 49088
rect 22428 49076 22434 49088
rect 24397 49079 24455 49085
rect 24397 49076 24409 49079
rect 22428 49048 24409 49076
rect 22428 49036 22434 49048
rect 24397 49045 24409 49048
rect 24443 49045 24455 49079
rect 24397 49039 24455 49045
rect 25406 49036 25412 49088
rect 25464 49076 25470 49088
rect 26053 49079 26111 49085
rect 26053 49076 26065 49079
rect 25464 49048 26065 49076
rect 25464 49036 25470 49048
rect 26053 49045 26065 49048
rect 26099 49045 26111 49079
rect 26053 49039 26111 49045
rect 32122 49036 32128 49088
rect 32180 49076 32186 49088
rect 32217 49079 32275 49085
rect 32217 49076 32229 49079
rect 32180 49048 32229 49076
rect 32180 49036 32186 49048
rect 32217 49045 32229 49048
rect 32263 49045 32275 49079
rect 32217 49039 32275 49045
rect 38010 49036 38016 49088
rect 38068 49076 38074 49088
rect 38289 49079 38347 49085
rect 38289 49076 38301 49079
rect 38068 49048 38301 49076
rect 38068 49036 38074 49048
rect 38289 49045 38301 49048
rect 38335 49045 38347 49079
rect 40862 49076 40868 49088
rect 40823 49048 40868 49076
rect 38289 49039 38347 49045
rect 40862 49036 40868 49048
rect 40920 49036 40926 49088
rect 41598 49076 41604 49088
rect 41559 49048 41604 49076
rect 41598 49036 41604 49048
rect 41656 49036 41662 49088
rect 47302 49036 47308 49088
rect 47360 49076 47366 49088
rect 47857 49079 47915 49085
rect 47857 49076 47869 49079
rect 47360 49048 47869 49076
rect 47360 49036 47366 49048
rect 47857 49045 47869 49048
rect 47903 49045 47915 49079
rect 47857 49039 47915 49045
rect 1104 48986 48852 49008
rect 1104 48934 19574 48986
rect 19626 48934 19638 48986
rect 19690 48934 19702 48986
rect 19754 48934 19766 48986
rect 19818 48934 19830 48986
rect 19882 48934 48852 48986
rect 1104 48912 48852 48934
rect 41782 48872 41788 48884
rect 41743 48844 41788 48872
rect 41782 48832 41788 48844
rect 41840 48832 41846 48884
rect 48314 48872 48320 48884
rect 44744 48844 48320 48872
rect 2866 48764 2872 48816
rect 2924 48804 2930 48816
rect 3513 48807 3571 48813
rect 3513 48804 3525 48807
rect 2924 48776 3525 48804
rect 2924 48764 2930 48776
rect 3513 48773 3525 48776
rect 3559 48773 3571 48807
rect 3513 48767 3571 48773
rect 5534 48764 5540 48816
rect 5592 48804 5598 48816
rect 9309 48807 9367 48813
rect 5592 48776 7788 48804
rect 5592 48764 5598 48776
rect 1673 48671 1731 48677
rect 1673 48637 1685 48671
rect 1719 48637 1731 48671
rect 1673 48631 1731 48637
rect 1857 48671 1915 48677
rect 1857 48637 1869 48671
rect 1903 48668 1915 48671
rect 3050 48668 3056 48680
rect 1903 48640 3056 48668
rect 1903 48637 1915 48640
rect 1857 48631 1915 48637
rect 1688 48532 1716 48631
rect 3050 48628 3056 48640
rect 3108 48628 3114 48680
rect 3973 48671 4031 48677
rect 3973 48637 3985 48671
rect 4019 48637 4031 48671
rect 3973 48631 4031 48637
rect 4157 48671 4215 48677
rect 4157 48637 4169 48671
rect 4203 48668 4215 48671
rect 4890 48668 4896 48680
rect 4203 48640 4896 48668
rect 4203 48637 4215 48640
rect 4157 48631 4215 48637
rect 3988 48600 4016 48631
rect 4890 48628 4896 48640
rect 4948 48628 4954 48680
rect 5626 48668 5632 48680
rect 5587 48640 5632 48668
rect 5626 48628 5632 48640
rect 5684 48628 5690 48680
rect 6362 48668 6368 48680
rect 6323 48640 6368 48668
rect 6362 48628 6368 48640
rect 6420 48628 6426 48680
rect 6549 48671 6607 48677
rect 6549 48637 6561 48671
rect 6595 48668 6607 48671
rect 7558 48668 7564 48680
rect 6595 48640 7564 48668
rect 6595 48637 6607 48640
rect 6549 48631 6607 48637
rect 7558 48628 7564 48640
rect 7616 48628 7622 48680
rect 7760 48677 7788 48776
rect 9309 48773 9321 48807
rect 9355 48804 9367 48807
rect 10502 48804 10508 48816
rect 9355 48776 10508 48804
rect 9355 48773 9367 48776
rect 9309 48767 9367 48773
rect 10502 48764 10508 48776
rect 10560 48764 10566 48816
rect 34790 48764 34796 48816
rect 34848 48804 34854 48816
rect 35069 48807 35127 48813
rect 35069 48804 35081 48807
rect 34848 48776 35081 48804
rect 34848 48764 34854 48776
rect 35069 48773 35081 48776
rect 35115 48773 35127 48807
rect 36722 48804 36728 48816
rect 36683 48776 36728 48804
rect 35069 48767 35127 48773
rect 36722 48764 36728 48776
rect 36780 48764 36786 48816
rect 44744 48813 44772 48844
rect 48314 48832 48320 48844
rect 48372 48832 48378 48884
rect 44729 48807 44787 48813
rect 44729 48773 44741 48807
rect 44775 48773 44787 48807
rect 47762 48804 47768 48816
rect 47723 48776 47768 48804
rect 44729 48767 44787 48773
rect 47762 48764 47768 48776
rect 47820 48764 47826 48816
rect 18046 48696 18052 48748
rect 18104 48736 18110 48748
rect 19153 48739 19211 48745
rect 19153 48736 19165 48739
rect 18104 48708 19165 48736
rect 18104 48696 18110 48708
rect 19153 48705 19165 48708
rect 19199 48705 19211 48739
rect 19153 48699 19211 48705
rect 21269 48739 21327 48745
rect 21269 48705 21281 48739
rect 21315 48736 21327 48739
rect 21818 48736 21824 48748
rect 21315 48708 21824 48736
rect 21315 48705 21327 48708
rect 21269 48699 21327 48705
rect 21818 48696 21824 48708
rect 21876 48696 21882 48748
rect 32122 48736 32128 48748
rect 32083 48708 32128 48736
rect 32122 48696 32128 48708
rect 32180 48696 32186 48748
rect 34882 48736 34888 48748
rect 34843 48708 34888 48736
rect 34882 48696 34888 48708
rect 34940 48696 34946 48748
rect 41690 48736 41696 48748
rect 41651 48708 41696 48736
rect 41690 48696 41696 48708
rect 41748 48696 41754 48748
rect 7745 48671 7803 48677
rect 7745 48637 7757 48671
rect 7791 48637 7803 48671
rect 9122 48668 9128 48680
rect 9083 48640 9128 48668
rect 7745 48631 7803 48637
rect 9122 48628 9128 48640
rect 9180 48628 9186 48680
rect 9674 48668 9680 48680
rect 9635 48640 9680 48668
rect 9674 48628 9680 48640
rect 9732 48628 9738 48680
rect 12434 48628 12440 48680
rect 12492 48668 12498 48680
rect 12621 48671 12679 48677
rect 12492 48640 12537 48668
rect 12492 48628 12498 48640
rect 12621 48637 12633 48671
rect 12667 48668 12679 48671
rect 12802 48668 12808 48680
rect 12667 48640 12808 48668
rect 12667 48637 12679 48640
rect 12621 48631 12679 48637
rect 12802 48628 12808 48640
rect 12860 48628 12866 48680
rect 12897 48671 12955 48677
rect 12897 48637 12909 48671
rect 12943 48637 12955 48671
rect 12897 48631 12955 48637
rect 16117 48671 16175 48677
rect 16117 48637 16129 48671
rect 16163 48668 16175 48671
rect 16669 48671 16727 48677
rect 16669 48668 16681 48671
rect 16163 48640 16681 48668
rect 16163 48637 16175 48640
rect 16117 48631 16175 48637
rect 16669 48637 16681 48640
rect 16715 48637 16727 48671
rect 16850 48668 16856 48680
rect 16811 48640 16856 48668
rect 16669 48631 16727 48637
rect 4706 48600 4712 48612
rect 3988 48572 4712 48600
rect 4706 48560 4712 48572
rect 4764 48560 4770 48612
rect 12526 48560 12532 48612
rect 12584 48600 12590 48612
rect 12912 48600 12940 48631
rect 16850 48628 16856 48640
rect 16908 48628 16914 48680
rect 17034 48628 17040 48680
rect 17092 48668 17098 48680
rect 17129 48671 17187 48677
rect 17129 48668 17141 48671
rect 17092 48640 17141 48668
rect 17092 48628 17098 48640
rect 17129 48637 17141 48640
rect 17175 48637 17187 48671
rect 17129 48631 17187 48637
rect 22005 48671 22063 48677
rect 22005 48637 22017 48671
rect 22051 48668 22063 48671
rect 22465 48671 22523 48677
rect 22465 48668 22477 48671
rect 22051 48640 22477 48668
rect 22051 48637 22063 48640
rect 22005 48631 22063 48637
rect 22465 48637 22477 48640
rect 22511 48637 22523 48671
rect 22646 48668 22652 48680
rect 22607 48640 22652 48668
rect 22465 48631 22523 48637
rect 22646 48628 22652 48640
rect 22704 48628 22710 48680
rect 23474 48668 23480 48680
rect 23435 48640 23480 48668
rect 23474 48628 23480 48640
rect 23532 48628 23538 48680
rect 26421 48671 26479 48677
rect 26421 48637 26433 48671
rect 26467 48668 26479 48671
rect 27065 48671 27123 48677
rect 27065 48668 27077 48671
rect 26467 48640 27077 48668
rect 26467 48637 26479 48640
rect 26421 48631 26479 48637
rect 27065 48637 27077 48640
rect 27111 48637 27123 48671
rect 27246 48668 27252 48680
rect 27207 48640 27252 48668
rect 27065 48631 27123 48637
rect 27246 48628 27252 48640
rect 27304 48628 27310 48680
rect 27798 48668 27804 48680
rect 27759 48640 27804 48668
rect 27798 48628 27804 48640
rect 27856 48628 27862 48680
rect 29270 48628 29276 48680
rect 29328 48668 29334 48680
rect 29365 48671 29423 48677
rect 29365 48668 29377 48671
rect 29328 48640 29377 48668
rect 29328 48628 29334 48640
rect 29365 48637 29377 48640
rect 29411 48637 29423 48671
rect 29546 48668 29552 48680
rect 29507 48640 29552 48668
rect 29365 48631 29423 48637
rect 29546 48628 29552 48640
rect 29604 48628 29610 48680
rect 29822 48668 29828 48680
rect 29783 48640 29828 48668
rect 29822 48628 29828 48640
rect 29880 48628 29886 48680
rect 32306 48668 32312 48680
rect 32267 48640 32312 48668
rect 32306 48628 32312 48640
rect 32364 48628 32370 48680
rect 33134 48668 33140 48680
rect 33095 48640 33140 48668
rect 33134 48628 33140 48640
rect 33192 48628 33198 48680
rect 38749 48671 38807 48677
rect 38749 48637 38761 48671
rect 38795 48668 38807 48671
rect 39209 48671 39267 48677
rect 39209 48668 39221 48671
rect 38795 48640 39221 48668
rect 38795 48637 38807 48640
rect 38749 48631 38807 48637
rect 39209 48637 39221 48640
rect 39255 48637 39267 48671
rect 39390 48668 39396 48680
rect 39351 48640 39396 48668
rect 39209 48631 39267 48637
rect 39390 48628 39396 48640
rect 39448 48628 39454 48680
rect 40034 48668 40040 48680
rect 39995 48640 40040 48668
rect 40034 48628 40040 48640
rect 40092 48628 40098 48680
rect 41414 48628 41420 48680
rect 41472 48668 41478 48680
rect 42889 48671 42947 48677
rect 42889 48668 42901 48671
rect 41472 48640 42901 48668
rect 41472 48628 41478 48640
rect 42889 48637 42901 48640
rect 42935 48637 42947 48671
rect 43070 48668 43076 48680
rect 43031 48640 43076 48668
rect 42889 48631 42947 48637
rect 43070 48628 43076 48640
rect 43128 48628 43134 48680
rect 44818 48628 44824 48680
rect 44876 48668 44882 48680
rect 45189 48671 45247 48677
rect 45189 48668 45201 48671
rect 44876 48640 45201 48668
rect 44876 48628 44882 48640
rect 45189 48637 45201 48640
rect 45235 48637 45247 48671
rect 45370 48668 45376 48680
rect 45331 48640 45376 48668
rect 45189 48631 45247 48637
rect 45370 48628 45376 48640
rect 45428 48628 45434 48680
rect 45738 48668 45744 48680
rect 45699 48640 45744 48668
rect 45738 48628 45744 48640
rect 45796 48628 45802 48680
rect 12584 48572 12940 48600
rect 12584 48560 12590 48572
rect 5350 48532 5356 48544
rect 1688 48504 5356 48532
rect 5350 48492 5356 48504
rect 5408 48492 5414 48544
rect 11698 48532 11704 48544
rect 11659 48504 11704 48532
rect 11698 48492 11704 48504
rect 11756 48492 11762 48544
rect 14918 48532 14924 48544
rect 14879 48504 14924 48532
rect 14918 48492 14924 48504
rect 14976 48492 14982 48544
rect 18046 48492 18052 48544
rect 18104 48532 18110 48544
rect 18969 48535 19027 48541
rect 18969 48532 18981 48535
rect 18104 48504 18981 48532
rect 18104 48492 18110 48504
rect 18969 48501 18981 48504
rect 19015 48501 19027 48535
rect 20438 48532 20444 48544
rect 20399 48504 20444 48532
rect 18969 48495 19027 48501
rect 20438 48492 20444 48504
rect 20496 48492 20502 48544
rect 24946 48532 24952 48544
rect 24907 48504 24952 48532
rect 24946 48492 24952 48504
rect 25004 48492 25010 48544
rect 25777 48535 25835 48541
rect 25777 48501 25789 48535
rect 25823 48532 25835 48535
rect 26694 48532 26700 48544
rect 25823 48504 26700 48532
rect 25823 48501 25835 48504
rect 25777 48495 25835 48501
rect 26694 48492 26700 48504
rect 26752 48492 26758 48544
rect 47118 48492 47124 48544
rect 47176 48532 47182 48544
rect 47857 48535 47915 48541
rect 47857 48532 47869 48535
rect 47176 48504 47869 48532
rect 47176 48492 47182 48504
rect 47857 48501 47869 48504
rect 47903 48501 47915 48535
rect 47857 48495 47915 48501
rect 1104 48442 48852 48464
rect 1104 48390 4214 48442
rect 4266 48390 4278 48442
rect 4330 48390 4342 48442
rect 4394 48390 4406 48442
rect 4458 48390 4470 48442
rect 4522 48390 34934 48442
rect 34986 48390 34998 48442
rect 35050 48390 35062 48442
rect 35114 48390 35126 48442
rect 35178 48390 35190 48442
rect 35242 48390 48852 48442
rect 1104 48368 48852 48390
rect 3418 48288 3424 48340
rect 3476 48328 3482 48340
rect 6638 48328 6644 48340
rect 3476 48300 6644 48328
rect 3476 48288 3482 48300
rect 6638 48288 6644 48300
rect 6696 48288 6702 48340
rect 12434 48288 12440 48340
rect 12492 48328 12498 48340
rect 12713 48331 12771 48337
rect 12713 48328 12725 48331
rect 12492 48300 12725 48328
rect 12492 48288 12498 48300
rect 12713 48297 12725 48300
rect 12759 48297 12771 48331
rect 12713 48291 12771 48297
rect 12802 48288 12808 48340
rect 12860 48328 12866 48340
rect 13449 48331 13507 48337
rect 13449 48328 13461 48331
rect 12860 48300 13461 48328
rect 12860 48288 12866 48300
rect 13449 48297 13461 48300
rect 13495 48297 13507 48331
rect 13449 48291 13507 48297
rect 22646 48288 22652 48340
rect 22704 48328 22710 48340
rect 22925 48331 22983 48337
rect 22925 48328 22937 48331
rect 22704 48300 22937 48328
rect 22704 48288 22710 48300
rect 22925 48297 22937 48300
rect 22971 48297 22983 48331
rect 22925 48291 22983 48297
rect 24412 48300 25176 48328
rect 14 48220 20 48272
rect 72 48260 78 48272
rect 2774 48260 2780 48272
rect 72 48232 2780 48260
rect 72 48220 78 48232
rect 2774 48220 2780 48232
rect 2832 48220 2838 48272
rect 3970 48220 3976 48272
rect 4028 48260 4034 48272
rect 7374 48260 7380 48272
rect 4028 48232 5672 48260
rect 7335 48232 7380 48260
rect 4028 48220 4034 48232
rect 1302 48152 1308 48204
rect 1360 48192 1366 48204
rect 1857 48195 1915 48201
rect 1857 48192 1869 48195
rect 1360 48164 1869 48192
rect 1360 48152 1366 48164
rect 1857 48161 1869 48164
rect 1903 48161 1915 48195
rect 1857 48155 1915 48161
rect 4525 48195 4583 48201
rect 4525 48161 4537 48195
rect 4571 48192 4583 48195
rect 5534 48192 5540 48204
rect 4571 48164 5540 48192
rect 4571 48161 4583 48164
rect 4525 48155 4583 48161
rect 5534 48152 5540 48164
rect 5592 48152 5598 48204
rect 5644 48201 5672 48232
rect 7374 48220 7380 48232
rect 7432 48220 7438 48272
rect 7558 48220 7564 48272
rect 7616 48260 7622 48272
rect 8021 48263 8079 48269
rect 8021 48260 8033 48263
rect 7616 48232 8033 48260
rect 7616 48220 7622 48232
rect 8021 48229 8033 48232
rect 8067 48229 8079 48263
rect 8021 48223 8079 48229
rect 17402 48220 17408 48272
rect 17460 48260 17466 48272
rect 24412 48260 24440 48300
rect 17460 48232 18092 48260
rect 17460 48220 17466 48232
rect 5629 48195 5687 48201
rect 5629 48161 5641 48195
rect 5675 48161 5687 48195
rect 5629 48155 5687 48161
rect 9122 48152 9128 48204
rect 9180 48192 9186 48204
rect 9217 48195 9275 48201
rect 9217 48192 9229 48195
rect 9180 48164 9229 48192
rect 9180 48152 9186 48164
rect 9217 48161 9229 48164
rect 9263 48161 9275 48195
rect 9217 48155 9275 48161
rect 9861 48195 9919 48201
rect 9861 48161 9873 48195
rect 9907 48192 9919 48195
rect 11698 48192 11704 48204
rect 9907 48164 11704 48192
rect 9907 48161 9919 48164
rect 9861 48155 9919 48161
rect 11698 48152 11704 48164
rect 11756 48152 11762 48204
rect 14461 48195 14519 48201
rect 14461 48161 14473 48195
rect 14507 48192 14519 48195
rect 14918 48192 14924 48204
rect 14507 48164 14924 48192
rect 14507 48161 14519 48164
rect 14461 48155 14519 48161
rect 14918 48152 14924 48164
rect 14976 48152 14982 48204
rect 15010 48152 15016 48204
rect 15068 48192 15074 48204
rect 15197 48195 15255 48201
rect 15197 48192 15209 48195
rect 15068 48164 15209 48192
rect 15068 48152 15074 48164
rect 15197 48161 15209 48164
rect 15243 48161 15255 48195
rect 15197 48155 15255 48161
rect 16853 48195 16911 48201
rect 16853 48161 16865 48195
rect 16899 48192 16911 48195
rect 17954 48192 17960 48204
rect 16899 48164 17960 48192
rect 16899 48161 16911 48164
rect 16853 48155 16911 48161
rect 17954 48152 17960 48164
rect 18012 48152 18018 48204
rect 18064 48201 18092 48232
rect 22848 48232 24440 48260
rect 18049 48195 18107 48201
rect 18049 48161 18061 48195
rect 18095 48161 18107 48195
rect 18049 48155 18107 48161
rect 20257 48195 20315 48201
rect 20257 48161 20269 48195
rect 20303 48192 20315 48195
rect 20438 48192 20444 48204
rect 20303 48164 20444 48192
rect 20303 48161 20315 48164
rect 20257 48155 20315 48161
rect 20438 48152 20444 48164
rect 20496 48152 20502 48204
rect 20622 48152 20628 48204
rect 20680 48192 20686 48204
rect 20717 48195 20775 48201
rect 20717 48192 20729 48195
rect 20680 48164 20729 48192
rect 20680 48152 20686 48164
rect 20717 48161 20729 48164
rect 20763 48161 20775 48195
rect 20717 48155 20775 48161
rect 1397 48127 1455 48133
rect 1397 48093 1409 48127
rect 1443 48093 1455 48127
rect 3786 48124 3792 48136
rect 3747 48096 3792 48124
rect 1397 48087 1455 48093
rect 1412 47988 1440 48087
rect 3786 48084 3792 48096
rect 3844 48084 3850 48136
rect 7190 48084 7196 48136
rect 7248 48124 7254 48136
rect 7285 48127 7343 48133
rect 7285 48124 7297 48127
rect 7248 48096 7297 48124
rect 7248 48084 7254 48096
rect 7285 48093 7297 48096
rect 7331 48093 7343 48127
rect 7926 48124 7932 48136
rect 7887 48096 7932 48124
rect 7285 48087 7343 48093
rect 7926 48084 7932 48096
rect 7984 48084 7990 48136
rect 22848 48133 22876 48232
rect 24486 48220 24492 48272
rect 24544 48260 24550 48272
rect 25148 48260 25176 48300
rect 29546 48288 29552 48340
rect 29604 48328 29610 48340
rect 29641 48331 29699 48337
rect 29641 48328 29653 48331
rect 29604 48300 29653 48328
rect 29604 48288 29610 48300
rect 29641 48297 29653 48300
rect 29687 48297 29699 48331
rect 34790 48328 34796 48340
rect 34751 48300 34796 48328
rect 29641 48291 29699 48297
rect 34790 48288 34796 48300
rect 34848 48288 34854 48340
rect 39390 48288 39396 48340
rect 39448 48328 39454 48340
rect 39945 48331 40003 48337
rect 39945 48328 39957 48331
rect 39448 48300 39957 48328
rect 39448 48288 39454 48300
rect 39945 48297 39957 48300
rect 39991 48297 40003 48331
rect 39945 48291 40003 48297
rect 30650 48260 30656 48272
rect 24544 48232 25084 48260
rect 25148 48232 29684 48260
rect 30611 48232 30656 48260
rect 24544 48220 24550 48232
rect 24397 48195 24455 48201
rect 24397 48161 24409 48195
rect 24443 48192 24455 48195
rect 24946 48192 24952 48204
rect 24443 48164 24952 48192
rect 24443 48161 24455 48164
rect 24397 48155 24455 48161
rect 24946 48152 24952 48164
rect 25004 48152 25010 48204
rect 25056 48201 25084 48232
rect 25041 48195 25099 48201
rect 25041 48161 25053 48195
rect 25087 48161 25099 48195
rect 26694 48192 26700 48204
rect 26655 48164 26700 48192
rect 25041 48155 25099 48161
rect 26694 48152 26700 48164
rect 26752 48152 26758 48204
rect 27062 48152 27068 48204
rect 27120 48192 27126 48204
rect 27157 48195 27215 48201
rect 27157 48192 27169 48195
rect 27120 48164 27169 48192
rect 27120 48152 27126 48164
rect 27157 48161 27169 48164
rect 27203 48161 27215 48195
rect 27157 48155 27215 48161
rect 13357 48127 13415 48133
rect 13357 48093 13369 48127
rect 13403 48093 13415 48127
rect 13357 48087 13415 48093
rect 22833 48127 22891 48133
rect 22833 48093 22845 48127
rect 22879 48093 22891 48127
rect 23658 48124 23664 48136
rect 23619 48096 23664 48124
rect 22833 48087 22891 48093
rect 1578 48056 1584 48068
rect 1539 48028 1584 48056
rect 1578 48016 1584 48028
rect 1636 48016 1642 48068
rect 4709 48059 4767 48065
rect 4709 48025 4721 48059
rect 4755 48056 4767 48059
rect 4982 48056 4988 48068
rect 4755 48028 4988 48056
rect 4755 48025 4767 48028
rect 4709 48019 4767 48025
rect 4982 48016 4988 48028
rect 5040 48016 5046 48068
rect 10042 48056 10048 48068
rect 10003 48028 10048 48056
rect 10042 48016 10048 48028
rect 10100 48016 10106 48068
rect 10318 48016 10324 48068
rect 10376 48056 10382 48068
rect 11701 48059 11759 48065
rect 11701 48056 11713 48059
rect 10376 48028 11713 48056
rect 10376 48016 10382 48028
rect 11701 48025 11713 48028
rect 11747 48025 11759 48059
rect 11701 48019 11759 48025
rect 3878 47988 3884 48000
rect 1412 47960 3884 47988
rect 3878 47948 3884 47960
rect 3936 47948 3942 48000
rect 3973 47991 4031 47997
rect 3973 47957 3985 47991
rect 4019 47988 4031 47991
rect 4062 47988 4068 48000
rect 4019 47960 4068 47988
rect 4019 47957 4031 47960
rect 3973 47951 4031 47957
rect 4062 47948 4068 47960
rect 4120 47948 4126 48000
rect 13372 47988 13400 48087
rect 23658 48084 23664 48096
rect 23716 48084 23722 48136
rect 29546 48124 29552 48136
rect 29507 48096 29552 48124
rect 29546 48084 29552 48096
rect 29604 48084 29610 48136
rect 29656 48124 29684 48232
rect 30650 48220 30656 48232
rect 30708 48220 30714 48272
rect 36630 48220 36636 48272
rect 36688 48260 36694 48272
rect 44085 48263 44143 48269
rect 44085 48260 44097 48263
rect 36688 48232 44097 48260
rect 36688 48220 36694 48232
rect 44085 48229 44097 48232
rect 44131 48229 44143 48263
rect 44085 48223 44143 48229
rect 47026 48220 47032 48272
rect 47084 48260 47090 48272
rect 49602 48260 49608 48272
rect 47084 48232 49608 48260
rect 47084 48220 47090 48232
rect 49602 48220 49608 48232
rect 49660 48220 49666 48272
rect 31297 48195 31355 48201
rect 31297 48161 31309 48195
rect 31343 48192 31355 48195
rect 31938 48192 31944 48204
rect 31343 48164 31944 48192
rect 31343 48161 31355 48164
rect 31297 48155 31355 48161
rect 31938 48152 31944 48164
rect 31996 48152 32002 48204
rect 32214 48192 32220 48204
rect 32175 48164 32220 48192
rect 32214 48152 32220 48164
rect 32272 48152 32278 48204
rect 35437 48195 35495 48201
rect 35437 48161 35449 48195
rect 35483 48192 35495 48195
rect 36170 48192 36176 48204
rect 35483 48164 36176 48192
rect 35483 48161 35495 48164
rect 35437 48155 35495 48161
rect 36170 48152 36176 48164
rect 36228 48152 36234 48204
rect 36262 48152 36268 48204
rect 36320 48192 36326 48204
rect 42518 48192 42524 48204
rect 36320 48164 36365 48192
rect 42479 48164 42524 48192
rect 36320 48152 36326 48164
rect 42518 48152 42524 48164
rect 42576 48152 42582 48204
rect 46293 48195 46351 48201
rect 46293 48161 46305 48195
rect 46339 48192 46351 48195
rect 46658 48192 46664 48204
rect 46339 48164 46664 48192
rect 46339 48161 46351 48164
rect 46293 48155 46351 48161
rect 46658 48152 46664 48164
rect 46716 48152 46722 48204
rect 46842 48192 46848 48204
rect 46803 48164 46848 48192
rect 46842 48152 46848 48164
rect 46900 48152 46906 48204
rect 30558 48124 30564 48136
rect 29656 48096 30564 48124
rect 30558 48084 30564 48096
rect 30616 48084 30622 48136
rect 33318 48124 33324 48136
rect 32692 48096 33324 48124
rect 14366 48016 14372 48068
rect 14424 48056 14430 48068
rect 14645 48059 14703 48065
rect 14645 48056 14657 48059
rect 14424 48028 14657 48056
rect 14424 48016 14430 48028
rect 14645 48025 14657 48028
rect 14691 48025 14703 48059
rect 14645 48019 14703 48025
rect 17037 48059 17095 48065
rect 17037 48025 17049 48059
rect 17083 48056 17095 48059
rect 17402 48056 17408 48068
rect 17083 48028 17408 48056
rect 17083 48025 17095 48028
rect 17037 48019 17095 48025
rect 17402 48016 17408 48028
rect 17460 48016 17466 48068
rect 20254 48016 20260 48068
rect 20312 48056 20318 48068
rect 20441 48059 20499 48065
rect 20441 48056 20453 48059
rect 20312 48028 20453 48056
rect 20312 48016 20318 48028
rect 20441 48025 20453 48028
rect 20487 48025 20499 48059
rect 23566 48056 23572 48068
rect 20441 48019 20499 48025
rect 22066 48028 23572 48056
rect 16666 47988 16672 48000
rect 13372 47960 16672 47988
rect 16666 47948 16672 47960
rect 16724 47948 16730 48000
rect 17126 47948 17132 48000
rect 17184 47988 17190 48000
rect 22066 47988 22094 48028
rect 23566 48016 23572 48028
rect 23624 48016 23630 48068
rect 23753 48059 23811 48065
rect 23753 48025 23765 48059
rect 23799 48056 23811 48059
rect 24581 48059 24639 48065
rect 24581 48056 24593 48059
rect 23799 48028 24593 48056
rect 23799 48025 23811 48028
rect 23753 48019 23811 48025
rect 24581 48025 24593 48028
rect 24627 48025 24639 48059
rect 24581 48019 24639 48025
rect 26326 48016 26332 48068
rect 26384 48056 26390 48068
rect 26881 48059 26939 48065
rect 26881 48056 26893 48059
rect 26384 48028 26893 48056
rect 26384 48016 26390 48028
rect 26881 48025 26893 48028
rect 26927 48025 26939 48059
rect 26881 48019 26939 48025
rect 31110 48016 31116 48068
rect 31168 48056 31174 48068
rect 31481 48059 31539 48065
rect 31481 48056 31493 48059
rect 31168 48028 31493 48056
rect 31168 48016 31174 48028
rect 31481 48025 31493 48028
rect 31527 48025 31539 48059
rect 31481 48019 31539 48025
rect 17184 47960 22094 47988
rect 17184 47948 17190 47960
rect 24026 47948 24032 48000
rect 24084 47988 24090 48000
rect 32692 47988 32720 48096
rect 33318 48084 33324 48096
rect 33376 48124 33382 48136
rect 33597 48127 33655 48133
rect 33597 48124 33609 48127
rect 33376 48096 33609 48124
rect 33376 48084 33382 48096
rect 33597 48093 33609 48096
rect 33643 48093 33655 48127
rect 33597 48087 33655 48093
rect 34606 48084 34612 48136
rect 34664 48124 34670 48136
rect 34701 48127 34759 48133
rect 34701 48124 34713 48127
rect 34664 48096 34713 48124
rect 34664 48084 34670 48096
rect 34701 48093 34713 48096
rect 34747 48093 34759 48127
rect 34701 48087 34759 48093
rect 39853 48127 39911 48133
rect 39853 48093 39865 48127
rect 39899 48093 39911 48127
rect 39853 48087 39911 48093
rect 40957 48127 41015 48133
rect 40957 48093 40969 48127
rect 41003 48124 41015 48127
rect 41417 48127 41475 48133
rect 41417 48124 41429 48127
rect 41003 48096 41429 48124
rect 41003 48093 41015 48096
rect 40957 48087 41015 48093
rect 41417 48093 41429 48096
rect 41463 48093 41475 48127
rect 43898 48124 43904 48136
rect 43859 48096 43904 48124
rect 41417 48087 41475 48093
rect 35621 48059 35679 48065
rect 35621 48025 35633 48059
rect 35667 48056 35679 48059
rect 35894 48056 35900 48068
rect 35667 48028 35900 48056
rect 35667 48025 35679 48028
rect 35621 48019 35679 48025
rect 35894 48016 35900 48028
rect 35952 48016 35958 48068
rect 33686 47988 33692 48000
rect 24084 47960 32720 47988
rect 33647 47960 33692 47988
rect 24084 47948 24090 47960
rect 33686 47948 33692 47960
rect 33744 47948 33750 48000
rect 39868 47988 39896 48087
rect 43898 48084 43904 48096
rect 43956 48084 43962 48136
rect 44450 48084 44456 48136
rect 44508 48124 44514 48136
rect 45005 48127 45063 48133
rect 45005 48124 45017 48127
rect 44508 48096 45017 48124
rect 44508 48084 44514 48096
rect 45005 48093 45017 48096
rect 45051 48093 45063 48127
rect 45005 48087 45063 48093
rect 41601 48059 41659 48065
rect 41601 48025 41613 48059
rect 41647 48056 41659 48059
rect 41782 48056 41788 48068
rect 41647 48028 41788 48056
rect 41647 48025 41659 48028
rect 41601 48019 41659 48025
rect 41782 48016 41788 48028
rect 41840 48016 41846 48068
rect 46474 48056 46480 48068
rect 46435 48028 46480 48056
rect 46474 48016 46480 48028
rect 46532 48016 46538 48068
rect 44358 47988 44364 48000
rect 39868 47960 44364 47988
rect 44358 47948 44364 47960
rect 44416 47948 44422 48000
rect 44910 47948 44916 48000
rect 44968 47988 44974 48000
rect 45189 47991 45247 47997
rect 45189 47988 45201 47991
rect 44968 47960 45201 47988
rect 44968 47948 44974 47960
rect 45189 47957 45201 47960
rect 45235 47957 45247 47991
rect 45189 47951 45247 47957
rect 1104 47898 48852 47920
rect 1104 47846 19574 47898
rect 19626 47846 19638 47898
rect 19690 47846 19702 47898
rect 19754 47846 19766 47898
rect 19818 47846 19830 47898
rect 19882 47846 48852 47898
rect 1104 47824 48852 47846
rect 1578 47744 1584 47796
rect 1636 47784 1642 47796
rect 4341 47787 4399 47793
rect 4341 47784 4353 47787
rect 1636 47756 4353 47784
rect 1636 47744 1642 47756
rect 4341 47753 4353 47756
rect 4387 47753 4399 47787
rect 4982 47784 4988 47796
rect 4943 47756 4988 47784
rect 4341 47747 4399 47753
rect 4982 47744 4988 47756
rect 5040 47744 5046 47796
rect 9861 47787 9919 47793
rect 9861 47753 9873 47787
rect 9907 47784 9919 47787
rect 10042 47784 10048 47796
rect 9907 47756 10048 47784
rect 9907 47753 9919 47756
rect 9861 47747 9919 47753
rect 10042 47744 10048 47756
rect 10100 47744 10106 47796
rect 10502 47784 10508 47796
rect 10463 47756 10508 47784
rect 10502 47744 10508 47756
rect 10560 47744 10566 47796
rect 14366 47784 14372 47796
rect 14327 47756 14372 47784
rect 14366 47744 14372 47756
rect 14424 47744 14430 47796
rect 16761 47787 16819 47793
rect 16761 47753 16773 47787
rect 16807 47784 16819 47787
rect 16850 47784 16856 47796
rect 16807 47756 16856 47784
rect 16807 47753 16819 47756
rect 16761 47747 16819 47753
rect 16850 47744 16856 47756
rect 16908 47744 16914 47796
rect 17402 47784 17408 47796
rect 17363 47756 17408 47784
rect 17402 47744 17408 47756
rect 17460 47744 17466 47796
rect 20254 47784 20260 47796
rect 20215 47756 20260 47784
rect 20254 47744 20260 47756
rect 20312 47744 20318 47796
rect 22278 47784 22284 47796
rect 22239 47756 22284 47784
rect 22278 47744 22284 47756
rect 22336 47744 22342 47796
rect 26326 47784 26332 47796
rect 26287 47756 26332 47784
rect 26326 47744 26332 47756
rect 26384 47744 26390 47796
rect 27246 47744 27252 47796
rect 27304 47784 27310 47796
rect 27433 47787 27491 47793
rect 27433 47784 27445 47787
rect 27304 47756 27445 47784
rect 27304 47744 27310 47756
rect 27433 47753 27445 47756
rect 27479 47753 27491 47787
rect 31110 47784 31116 47796
rect 31071 47756 31116 47784
rect 27433 47747 27491 47753
rect 31110 47744 31116 47756
rect 31168 47744 31174 47796
rect 32306 47744 32312 47796
rect 32364 47784 32370 47796
rect 32493 47787 32551 47793
rect 32493 47784 32505 47787
rect 32364 47756 32505 47784
rect 32364 47744 32370 47756
rect 32493 47753 32505 47756
rect 32539 47753 32551 47787
rect 41690 47784 41696 47796
rect 32493 47747 32551 47753
rect 32600 47756 41696 47784
rect 5629 47719 5687 47725
rect 5629 47685 5641 47719
rect 5675 47716 5687 47719
rect 6178 47716 6184 47728
rect 5675 47688 6184 47716
rect 5675 47685 5687 47688
rect 5629 47679 5687 47685
rect 6178 47676 6184 47688
rect 6236 47676 6242 47728
rect 9784 47688 20852 47716
rect 4249 47651 4307 47657
rect 4249 47617 4261 47651
rect 4295 47648 4307 47651
rect 4798 47648 4804 47660
rect 4295 47620 4804 47648
rect 4295 47617 4307 47620
rect 4249 47611 4307 47617
rect 4798 47608 4804 47620
rect 4856 47608 4862 47660
rect 4893 47651 4951 47657
rect 4893 47617 4905 47651
rect 4939 47648 4951 47651
rect 6086 47648 6092 47660
rect 4939 47620 6092 47648
rect 4939 47617 4951 47620
rect 4893 47611 4951 47617
rect 6086 47608 6092 47620
rect 6144 47608 6150 47660
rect 8849 47651 8907 47657
rect 8849 47617 8861 47651
rect 8895 47648 8907 47651
rect 8938 47648 8944 47660
rect 8895 47620 8944 47648
rect 8895 47617 8907 47620
rect 8849 47611 8907 47617
rect 8938 47608 8944 47620
rect 8996 47608 9002 47660
rect 9784 47657 9812 47688
rect 9769 47651 9827 47657
rect 9769 47617 9781 47651
rect 9815 47617 9827 47651
rect 9769 47611 9827 47617
rect 10413 47651 10471 47657
rect 10413 47617 10425 47651
rect 10459 47648 10471 47651
rect 14274 47648 14280 47660
rect 10459 47620 14280 47648
rect 10459 47617 10471 47620
rect 10413 47611 10471 47617
rect 14274 47608 14280 47620
rect 14332 47608 14338 47660
rect 16666 47648 16672 47660
rect 16627 47620 16672 47648
rect 16666 47608 16672 47620
rect 16724 47608 16730 47660
rect 17313 47651 17371 47657
rect 17313 47617 17325 47651
rect 17359 47648 17371 47651
rect 17770 47648 17776 47660
rect 17359 47620 17776 47648
rect 17359 47617 17371 47620
rect 17313 47611 17371 47617
rect 17770 47608 17776 47620
rect 17828 47608 17834 47660
rect 20162 47648 20168 47660
rect 20123 47620 20168 47648
rect 20162 47608 20168 47620
rect 20220 47608 20226 47660
rect 20824 47657 20852 47688
rect 23566 47676 23572 47728
rect 23624 47716 23630 47728
rect 26510 47716 26516 47728
rect 23624 47688 26516 47716
rect 23624 47676 23630 47688
rect 20809 47651 20867 47657
rect 20809 47617 20821 47651
rect 20855 47648 20867 47651
rect 20990 47648 20996 47660
rect 20855 47620 20996 47648
rect 20855 47617 20867 47620
rect 20809 47611 20867 47617
rect 20990 47608 20996 47620
rect 21048 47608 21054 47660
rect 22189 47651 22247 47657
rect 22189 47617 22201 47651
rect 22235 47648 22247 47651
rect 22554 47648 22560 47660
rect 22235 47620 22560 47648
rect 22235 47617 22247 47620
rect 22189 47611 22247 47617
rect 22554 47608 22560 47620
rect 22612 47608 22618 47660
rect 26252 47657 26280 47688
rect 26510 47676 26516 47688
rect 26568 47716 26574 47728
rect 32600 47716 32628 47756
rect 41690 47744 41696 47756
rect 41748 47744 41754 47796
rect 41785 47787 41843 47793
rect 41785 47753 41797 47787
rect 41831 47784 41843 47787
rect 43070 47784 43076 47796
rect 41831 47756 43076 47784
rect 41831 47753 41843 47756
rect 41785 47747 41843 47753
rect 43070 47744 43076 47756
rect 43128 47744 43134 47796
rect 33686 47716 33692 47728
rect 26568 47688 32628 47716
rect 33647 47688 33692 47716
rect 26568 47676 26574 47688
rect 33686 47676 33692 47688
rect 33744 47676 33750 47728
rect 35894 47676 35900 47728
rect 35952 47716 35958 47728
rect 35952 47688 35997 47716
rect 35952 47676 35958 47688
rect 26237 47651 26295 47657
rect 26237 47617 26249 47651
rect 26283 47617 26295 47651
rect 26237 47611 26295 47617
rect 27154 47608 27160 47660
rect 27212 47648 27218 47660
rect 27341 47651 27399 47657
rect 27341 47648 27353 47651
rect 27212 47620 27353 47648
rect 27212 47608 27218 47620
rect 27341 47617 27353 47620
rect 27387 47617 27399 47651
rect 27982 47648 27988 47660
rect 27943 47620 27988 47648
rect 27341 47611 27399 47617
rect 27982 47608 27988 47620
rect 28040 47608 28046 47660
rect 30466 47648 30472 47660
rect 30427 47620 30472 47648
rect 30466 47608 30472 47620
rect 30524 47608 30530 47660
rect 31018 47648 31024 47660
rect 30979 47620 31024 47648
rect 31018 47608 31024 47620
rect 31076 47608 31082 47660
rect 32398 47648 32404 47660
rect 32359 47620 32404 47648
rect 32398 47608 32404 47620
rect 32456 47608 32462 47660
rect 33502 47648 33508 47660
rect 33463 47620 33508 47648
rect 33502 47608 33508 47620
rect 33560 47608 33566 47660
rect 35802 47648 35808 47660
rect 35763 47620 35808 47648
rect 35802 47608 35808 47620
rect 35860 47608 35866 47660
rect 41233 47651 41291 47657
rect 41233 47617 41245 47651
rect 41279 47648 41291 47651
rect 41414 47648 41420 47660
rect 41279 47620 41420 47648
rect 41279 47617 41291 47620
rect 41233 47611 41291 47617
rect 41414 47608 41420 47620
rect 41472 47608 41478 47660
rect 41708 47657 41736 47744
rect 43901 47719 43959 47725
rect 43901 47685 43913 47719
rect 43947 47716 43959 47719
rect 45554 47716 45560 47728
rect 43947 47688 45560 47716
rect 43947 47685 43959 47688
rect 43901 47679 43959 47685
rect 45554 47676 45560 47688
rect 45612 47676 45618 47728
rect 47762 47716 47768 47728
rect 47723 47688 47768 47716
rect 47762 47676 47768 47688
rect 47820 47676 47826 47728
rect 41693 47651 41751 47657
rect 41693 47617 41705 47651
rect 41739 47617 41751 47651
rect 41693 47611 41751 47617
rect 42521 47651 42579 47657
rect 42521 47617 42533 47651
rect 42567 47648 42579 47651
rect 42702 47648 42708 47660
rect 42567 47620 42708 47648
rect 42567 47617 42579 47620
rect 42521 47611 42579 47617
rect 1946 47580 1952 47592
rect 1907 47552 1952 47580
rect 1946 47540 1952 47552
rect 2004 47540 2010 47592
rect 2133 47583 2191 47589
rect 2133 47549 2145 47583
rect 2179 47580 2191 47583
rect 2866 47580 2872 47592
rect 2179 47552 2872 47580
rect 2179 47549 2191 47552
rect 2133 47543 2191 47549
rect 2866 47540 2872 47552
rect 2924 47540 2930 47592
rect 3142 47580 3148 47592
rect 3103 47552 3148 47580
rect 3142 47540 3148 47552
rect 3200 47540 3206 47592
rect 6365 47583 6423 47589
rect 6365 47549 6377 47583
rect 6411 47549 6423 47583
rect 6546 47580 6552 47592
rect 6507 47552 6552 47580
rect 6365 47543 6423 47549
rect 6380 47512 6408 47543
rect 6546 47540 6552 47552
rect 6604 47540 6610 47592
rect 6638 47540 6644 47592
rect 6696 47580 6702 47592
rect 6917 47583 6975 47589
rect 6917 47580 6929 47583
rect 6696 47552 6929 47580
rect 6696 47540 6702 47552
rect 6917 47549 6929 47552
rect 6963 47549 6975 47583
rect 26418 47580 26424 47592
rect 6917 47543 6975 47549
rect 9646 47552 26424 47580
rect 9646 47512 9674 47552
rect 26418 47540 26424 47552
rect 26476 47540 26482 47592
rect 28166 47580 28172 47592
rect 28127 47552 28172 47580
rect 28166 47540 28172 47552
rect 28224 47540 28230 47592
rect 28442 47580 28448 47592
rect 28403 47552 28448 47580
rect 28442 47540 28448 47552
rect 28500 47540 28506 47592
rect 34698 47580 34704 47592
rect 34659 47552 34704 47580
rect 34698 47540 34704 47552
rect 34756 47540 34762 47592
rect 41708 47580 41736 47611
rect 42702 47608 42708 47620
rect 42760 47648 42766 47660
rect 43625 47651 43683 47657
rect 43625 47648 43637 47651
rect 42760 47620 43637 47648
rect 42760 47608 42766 47620
rect 43625 47617 43637 47620
rect 43671 47617 43683 47651
rect 43625 47611 43683 47617
rect 42794 47580 42800 47592
rect 41708 47552 42800 47580
rect 42794 47540 42800 47552
rect 42852 47540 42858 47592
rect 43073 47583 43131 47589
rect 43073 47549 43085 47583
rect 43119 47549 43131 47583
rect 45094 47580 45100 47592
rect 45055 47552 45100 47580
rect 43073 47543 43131 47549
rect 6380 47484 9674 47512
rect 17402 47472 17408 47524
rect 17460 47512 17466 47524
rect 34606 47512 34612 47524
rect 17460 47484 34612 47512
rect 17460 47472 17466 47484
rect 34606 47472 34612 47484
rect 34664 47472 34670 47524
rect 5721 47447 5779 47453
rect 5721 47413 5733 47447
rect 5767 47444 5779 47447
rect 6638 47444 6644 47456
rect 5767 47416 6644 47444
rect 5767 47413 5779 47416
rect 5721 47407 5779 47413
rect 6638 47404 6644 47416
rect 6696 47404 6702 47456
rect 20530 47404 20536 47456
rect 20588 47444 20594 47456
rect 20901 47447 20959 47453
rect 20901 47444 20913 47447
rect 20588 47416 20913 47444
rect 20588 47404 20594 47416
rect 20901 47413 20913 47416
rect 20947 47413 20959 47447
rect 20901 47407 20959 47413
rect 20990 47404 20996 47456
rect 21048 47444 21054 47456
rect 31018 47444 31024 47456
rect 21048 47416 31024 47444
rect 21048 47404 21054 47416
rect 31018 47404 31024 47416
rect 31076 47444 31082 47456
rect 31294 47444 31300 47456
rect 31076 47416 31300 47444
rect 31076 47404 31082 47416
rect 31294 47404 31300 47416
rect 31352 47404 31358 47456
rect 43088 47444 43116 47543
rect 45094 47540 45100 47552
rect 45152 47540 45158 47592
rect 45278 47580 45284 47592
rect 45239 47552 45284 47580
rect 45278 47540 45284 47552
rect 45336 47540 45342 47592
rect 46566 47580 46572 47592
rect 46527 47552 46572 47580
rect 46566 47540 46572 47552
rect 46624 47540 46630 47592
rect 46566 47444 46572 47456
rect 43088 47416 46572 47444
rect 46566 47404 46572 47416
rect 46624 47404 46630 47456
rect 47578 47404 47584 47456
rect 47636 47444 47642 47456
rect 47857 47447 47915 47453
rect 47857 47444 47869 47447
rect 47636 47416 47869 47444
rect 47636 47404 47642 47416
rect 47857 47413 47869 47416
rect 47903 47413 47915 47447
rect 47857 47407 47915 47413
rect 1104 47354 48852 47376
rect 1104 47302 4214 47354
rect 4266 47302 4278 47354
rect 4330 47302 4342 47354
rect 4394 47302 4406 47354
rect 4458 47302 4470 47354
rect 4522 47302 34934 47354
rect 34986 47302 34998 47354
rect 35050 47302 35062 47354
rect 35114 47302 35126 47354
rect 35178 47302 35190 47354
rect 35242 47302 48852 47354
rect 1104 47280 48852 47302
rect 3050 47200 3056 47252
rect 3108 47240 3114 47252
rect 3881 47243 3939 47249
rect 3881 47240 3893 47243
rect 3108 47212 3893 47240
rect 3108 47200 3114 47212
rect 3881 47209 3893 47212
rect 3927 47209 3939 47243
rect 3881 47203 3939 47209
rect 4801 47243 4859 47249
rect 4801 47209 4813 47243
rect 4847 47240 4859 47243
rect 4890 47240 4896 47252
rect 4847 47212 4896 47240
rect 4847 47209 4859 47212
rect 4801 47203 4859 47209
rect 4890 47200 4896 47212
rect 4948 47200 4954 47252
rect 5534 47240 5540 47252
rect 5495 47212 5540 47240
rect 5534 47200 5540 47212
rect 5592 47200 5598 47252
rect 6273 47243 6331 47249
rect 6273 47209 6285 47243
rect 6319 47240 6331 47243
rect 6546 47240 6552 47252
rect 6319 47212 6552 47240
rect 6319 47209 6331 47212
rect 6273 47203 6331 47209
rect 6546 47200 6552 47212
rect 6604 47200 6610 47252
rect 6914 47200 6920 47252
rect 6972 47240 6978 47252
rect 7009 47243 7067 47249
rect 7009 47240 7021 47243
rect 6972 47212 7021 47240
rect 6972 47200 6978 47212
rect 7009 47209 7021 47212
rect 7055 47209 7067 47243
rect 7009 47203 7067 47209
rect 7837 47243 7895 47249
rect 7837 47209 7849 47243
rect 7883 47240 7895 47243
rect 8478 47240 8484 47252
rect 7883 47212 8484 47240
rect 7883 47209 7895 47212
rect 7837 47203 7895 47209
rect 8478 47200 8484 47212
rect 8536 47200 8542 47252
rect 10962 47200 10968 47252
rect 11020 47240 11026 47252
rect 13262 47240 13268 47252
rect 11020 47212 13268 47240
rect 11020 47200 11026 47212
rect 13262 47200 13268 47212
rect 13320 47200 13326 47252
rect 14274 47200 14280 47252
rect 14332 47240 14338 47252
rect 24026 47240 24032 47252
rect 14332 47212 24032 47240
rect 14332 47200 14338 47212
rect 24026 47200 24032 47212
rect 24084 47200 24090 47252
rect 27893 47243 27951 47249
rect 27893 47209 27905 47243
rect 27939 47240 27951 47243
rect 28166 47240 28172 47252
rect 27939 47212 28172 47240
rect 27939 47209 27951 47212
rect 27893 47203 27951 47209
rect 28166 47200 28172 47212
rect 28224 47200 28230 47252
rect 42334 47240 42340 47252
rect 31726 47212 42340 47240
rect 3602 47172 3608 47184
rect 1412 47144 3608 47172
rect 1412 47113 1440 47144
rect 3602 47132 3608 47144
rect 3660 47132 3666 47184
rect 17126 47172 17132 47184
rect 6886 47144 17132 47172
rect 1397 47107 1455 47113
rect 1397 47073 1409 47107
rect 1443 47073 1455 47107
rect 1854 47104 1860 47116
rect 1815 47076 1860 47104
rect 1397 47067 1455 47073
rect 1854 47064 1860 47076
rect 1912 47064 1918 47116
rect 6886 47104 6914 47144
rect 17126 47132 17132 47144
rect 17184 47132 17190 47184
rect 29546 47172 29552 47184
rect 17236 47144 20668 47172
rect 4724 47076 6914 47104
rect 3326 46996 3332 47048
rect 3384 47036 3390 47048
rect 4724 47045 4752 47076
rect 3789 47039 3847 47045
rect 3789 47036 3801 47039
rect 3384 47008 3801 47036
rect 3384 46996 3390 47008
rect 3789 47005 3801 47008
rect 3835 47005 3847 47039
rect 3789 46999 3847 47005
rect 4709 47039 4767 47045
rect 4709 47005 4721 47039
rect 4755 47005 4767 47039
rect 4709 46999 4767 47005
rect 6086 46996 6092 47048
rect 6144 47036 6150 47048
rect 6181 47039 6239 47045
rect 6181 47036 6193 47039
rect 6144 47008 6193 47036
rect 6144 46996 6150 47008
rect 6181 47005 6193 47008
rect 6227 47036 6239 47039
rect 7742 47036 7748 47048
rect 6227 47008 6914 47036
rect 7703 47008 7748 47036
rect 6227 47005 6239 47008
rect 6181 46999 6239 47005
rect 1578 46968 1584 46980
rect 1539 46940 1584 46968
rect 1578 46928 1584 46940
rect 1636 46928 1642 46980
rect 6886 46968 6914 47008
rect 7742 46996 7748 47008
rect 7800 46996 7806 47048
rect 7926 46996 7932 47048
rect 7984 47036 7990 47048
rect 17236 47036 17264 47144
rect 20530 47104 20536 47116
rect 20491 47076 20536 47104
rect 20530 47064 20536 47076
rect 20588 47064 20594 47116
rect 20640 47104 20668 47144
rect 20824 47144 29552 47172
rect 20824 47104 20852 47144
rect 29546 47132 29552 47144
rect 29604 47172 29610 47184
rect 31726 47172 31754 47212
rect 42334 47200 42340 47212
rect 42392 47200 42398 47252
rect 45097 47243 45155 47249
rect 45097 47209 45109 47243
rect 45143 47240 45155 47243
rect 45278 47240 45284 47252
rect 45143 47212 45284 47240
rect 45143 47209 45155 47212
rect 45097 47203 45155 47209
rect 45278 47200 45284 47212
rect 45336 47200 45342 47252
rect 29604 47144 31754 47172
rect 29604 47132 29610 47144
rect 35802 47132 35808 47184
rect 35860 47172 35866 47184
rect 35860 47144 41414 47172
rect 35860 47132 35866 47144
rect 32398 47104 32404 47116
rect 20640 47076 20852 47104
rect 22204 47076 32404 47104
rect 20346 47036 20352 47048
rect 7984 47008 17264 47036
rect 20307 47008 20352 47036
rect 7984 46996 7990 47008
rect 20346 46996 20352 47008
rect 20404 46996 20410 47048
rect 22204 47036 22232 47076
rect 32398 47064 32404 47076
rect 32456 47104 32462 47116
rect 33226 47104 33232 47116
rect 32456 47076 33232 47104
rect 32456 47064 32462 47076
rect 33226 47064 33232 47076
rect 33284 47064 33290 47116
rect 41386 47104 41414 47144
rect 43622 47104 43628 47116
rect 41386 47076 43628 47104
rect 43622 47064 43628 47076
rect 43680 47064 43686 47116
rect 44726 47064 44732 47116
rect 44784 47104 44790 47116
rect 46293 47107 46351 47113
rect 46293 47104 46305 47107
rect 44784 47076 46305 47104
rect 44784 47064 44790 47076
rect 46293 47073 46305 47076
rect 46339 47073 46351 47107
rect 46750 47104 46756 47116
rect 46711 47076 46756 47104
rect 46293 47067 46351 47073
rect 46750 47064 46756 47076
rect 46808 47064 46814 47116
rect 22066 47008 22232 47036
rect 27801 47039 27859 47045
rect 22066 46968 22094 47008
rect 27801 47005 27813 47039
rect 27847 47036 27859 47039
rect 28258 47036 28264 47048
rect 27847 47008 28264 47036
rect 27847 47005 27859 47008
rect 27801 46999 27859 47005
rect 28258 46996 28264 47008
rect 28316 46996 28322 47048
rect 41601 47039 41659 47045
rect 41601 47005 41613 47039
rect 41647 47036 41659 47039
rect 42702 47036 42708 47048
rect 41647 47008 42708 47036
rect 41647 47005 41659 47008
rect 41601 46999 41659 47005
rect 42702 46996 42708 47008
rect 42760 47036 42766 47048
rect 43257 47039 43315 47045
rect 43257 47036 43269 47039
rect 42760 47008 43269 47036
rect 42760 46996 42766 47008
rect 43257 47005 43269 47008
rect 43303 47005 43315 47039
rect 45002 47036 45008 47048
rect 44963 47008 45008 47036
rect 43257 46999 43315 47005
rect 45002 46996 45008 47008
rect 45060 46996 45066 47048
rect 45646 47036 45652 47048
rect 45607 47008 45652 47036
rect 45646 46996 45652 47008
rect 45704 46996 45710 47048
rect 47946 46996 47952 47048
rect 48004 47036 48010 47048
rect 48958 47036 48964 47048
rect 48004 47008 48964 47036
rect 48004 46996 48010 47008
rect 48958 46996 48964 47008
rect 49016 46996 49022 47048
rect 6886 46940 20300 46968
rect 20272 46939 20300 46940
rect 20456 46940 22094 46968
rect 22189 46971 22247 46977
rect 20456 46939 20484 46940
rect 20272 46911 20484 46939
rect 22189 46937 22201 46971
rect 22235 46968 22247 46971
rect 39298 46968 39304 46980
rect 22235 46940 39304 46968
rect 22235 46937 22247 46940
rect 22189 46931 22247 46937
rect 39298 46928 39304 46940
rect 39356 46928 39362 46980
rect 41506 46928 41512 46980
rect 41564 46968 41570 46980
rect 41782 46968 41788 46980
rect 41564 46940 41788 46968
rect 41564 46928 41570 46940
rect 41782 46928 41788 46940
rect 41840 46928 41846 46980
rect 42334 46968 42340 46980
rect 42295 46940 42340 46968
rect 42334 46928 42340 46940
rect 42392 46928 42398 46980
rect 45830 46928 45836 46980
rect 45888 46968 45894 46980
rect 46477 46971 46535 46977
rect 46477 46968 46489 46971
rect 45888 46940 46489 46968
rect 45888 46928 45894 46940
rect 46477 46937 46489 46940
rect 46523 46937 46535 46971
rect 46477 46931 46535 46937
rect 45738 46900 45744 46912
rect 45699 46872 45744 46900
rect 45738 46860 45744 46872
rect 45796 46860 45802 46912
rect 1104 46810 48852 46832
rect 1104 46758 19574 46810
rect 19626 46758 19638 46810
rect 19690 46758 19702 46810
rect 19754 46758 19766 46810
rect 19818 46758 19830 46810
rect 19882 46758 48852 46810
rect 1104 46736 48852 46758
rect 2866 46696 2872 46708
rect 2827 46668 2872 46696
rect 2866 46656 2872 46668
rect 2924 46656 2930 46708
rect 44082 46696 44088 46708
rect 44043 46668 44088 46696
rect 44082 46656 44088 46668
rect 44140 46656 44146 46708
rect 11514 46628 11520 46640
rect 2792 46600 11520 46628
rect 1581 46563 1639 46569
rect 1581 46529 1593 46563
rect 1627 46560 1639 46563
rect 1946 46560 1952 46572
rect 1627 46532 1952 46560
rect 1627 46529 1639 46532
rect 1581 46523 1639 46529
rect 1946 46520 1952 46532
rect 2004 46520 2010 46572
rect 2038 46520 2044 46572
rect 2096 46560 2102 46572
rect 2096 46532 2141 46560
rect 2096 46520 2102 46532
rect 2314 46520 2320 46572
rect 2372 46560 2378 46572
rect 2792 46569 2820 46600
rect 11514 46588 11520 46600
rect 11572 46588 11578 46640
rect 23658 46588 23664 46640
rect 23716 46628 23722 46640
rect 24762 46628 24768 46640
rect 23716 46600 24768 46628
rect 23716 46588 23722 46600
rect 24762 46588 24768 46600
rect 24820 46628 24826 46640
rect 45002 46628 45008 46640
rect 24820 46600 45008 46628
rect 24820 46588 24826 46600
rect 2777 46563 2835 46569
rect 2777 46560 2789 46563
rect 2372 46532 2789 46560
rect 2372 46520 2378 46532
rect 2777 46529 2789 46532
rect 2823 46529 2835 46563
rect 3602 46560 3608 46572
rect 3563 46532 3608 46560
rect 2777 46523 2835 46529
rect 3602 46520 3608 46532
rect 3660 46520 3666 46572
rect 4249 46563 4307 46569
rect 4249 46529 4261 46563
rect 4295 46560 4307 46563
rect 4706 46560 4712 46572
rect 4295 46532 4712 46560
rect 4295 46529 4307 46532
rect 4249 46523 4307 46529
rect 4706 46520 4712 46532
rect 4764 46520 4770 46572
rect 5350 46560 5356 46572
rect 5311 46532 5356 46560
rect 5350 46520 5356 46532
rect 5408 46520 5414 46572
rect 42613 46563 42671 46569
rect 42613 46529 42625 46563
rect 42659 46560 42671 46563
rect 42702 46560 42708 46572
rect 42659 46532 42708 46560
rect 42659 46529 42671 46532
rect 42613 46523 42671 46529
rect 42702 46520 42708 46532
rect 42760 46520 42766 46572
rect 44008 46569 44036 46600
rect 45002 46588 45008 46600
rect 45060 46588 45066 46640
rect 45373 46631 45431 46637
rect 45373 46597 45385 46631
rect 45419 46628 45431 46631
rect 45738 46628 45744 46640
rect 45419 46600 45744 46628
rect 45419 46597 45431 46600
rect 45373 46591 45431 46597
rect 45738 46588 45744 46600
rect 45796 46588 45802 46640
rect 47026 46628 47032 46640
rect 46987 46600 47032 46628
rect 47026 46588 47032 46600
rect 47084 46588 47090 46640
rect 47946 46628 47952 46640
rect 47907 46600 47952 46628
rect 47946 46588 47952 46600
rect 48004 46588 48010 46640
rect 43993 46563 44051 46569
rect 43993 46529 44005 46563
rect 44039 46529 44051 46563
rect 43993 46523 44051 46529
rect 42794 46492 42800 46504
rect 42755 46464 42800 46492
rect 42794 46452 42800 46464
rect 42852 46452 42858 46504
rect 44174 46452 44180 46504
rect 44232 46492 44238 46504
rect 45189 46495 45247 46501
rect 45189 46492 45201 46495
rect 44232 46464 45201 46492
rect 44232 46452 44238 46464
rect 45189 46461 45201 46464
rect 45235 46461 45247 46495
rect 45189 46455 45247 46461
rect 1762 46316 1768 46368
rect 1820 46356 1826 46368
rect 2225 46359 2283 46365
rect 2225 46356 2237 46359
rect 1820 46328 2237 46356
rect 1820 46316 1826 46328
rect 2225 46325 2237 46328
rect 2271 46325 2283 46359
rect 2225 46319 2283 46325
rect 47762 46316 47768 46368
rect 47820 46356 47826 46368
rect 48041 46359 48099 46365
rect 48041 46356 48053 46359
rect 47820 46328 48053 46356
rect 47820 46316 47826 46328
rect 48041 46325 48053 46328
rect 48087 46325 48099 46359
rect 48041 46319 48099 46325
rect 1104 46266 48852 46288
rect 1104 46214 4214 46266
rect 4266 46214 4278 46266
rect 4330 46214 4342 46266
rect 4394 46214 4406 46266
rect 4458 46214 4470 46266
rect 4522 46214 34934 46266
rect 34986 46214 34998 46266
rect 35050 46214 35062 46266
rect 35114 46214 35126 46266
rect 35178 46214 35190 46266
rect 35242 46214 48852 46266
rect 1104 46192 48852 46214
rect 1578 46112 1584 46164
rect 1636 46152 1642 46164
rect 2409 46155 2467 46161
rect 2409 46152 2421 46155
rect 1636 46124 2421 46152
rect 1636 46112 1642 46124
rect 2409 46121 2421 46124
rect 2455 46121 2467 46155
rect 2409 46115 2467 46121
rect 3878 46112 3884 46164
rect 3936 46152 3942 46164
rect 3973 46155 4031 46161
rect 3973 46152 3985 46155
rect 3936 46124 3985 46152
rect 3936 46112 3942 46124
rect 3973 46121 3985 46124
rect 4019 46121 4031 46155
rect 3973 46115 4031 46121
rect 42429 46155 42487 46161
rect 42429 46121 42441 46155
rect 42475 46152 42487 46155
rect 42702 46152 42708 46164
rect 42475 46124 42708 46152
rect 42475 46121 42487 46124
rect 42429 46115 42487 46121
rect 42702 46112 42708 46124
rect 42760 46112 42766 46164
rect 43809 46155 43867 46161
rect 43809 46121 43821 46155
rect 43855 46152 43867 46155
rect 43990 46152 43996 46164
rect 43855 46124 43996 46152
rect 43855 46121 43867 46124
rect 43809 46115 43867 46121
rect 43990 46112 43996 46124
rect 44048 46112 44054 46164
rect 44453 46155 44511 46161
rect 44453 46121 44465 46155
rect 44499 46152 44511 46155
rect 44818 46152 44824 46164
rect 44499 46124 44824 46152
rect 44499 46121 44511 46124
rect 44453 46115 44511 46121
rect 44818 46112 44824 46124
rect 44876 46112 44882 46164
rect 45097 46155 45155 46161
rect 45097 46121 45109 46155
rect 45143 46152 45155 46155
rect 45370 46152 45376 46164
rect 45143 46124 45376 46152
rect 45143 46121 45155 46124
rect 45097 46115 45155 46121
rect 45370 46112 45376 46124
rect 45428 46112 45434 46164
rect 45741 46155 45799 46161
rect 45741 46121 45753 46155
rect 45787 46152 45799 46155
rect 46474 46152 46480 46164
rect 45787 46124 46480 46152
rect 45787 46121 45799 46124
rect 45741 46115 45799 46121
rect 46474 46112 46480 46124
rect 46532 46112 46538 46164
rect 30558 46044 30564 46096
rect 30616 46084 30622 46096
rect 31662 46084 31668 46096
rect 30616 46056 31668 46084
rect 30616 46044 30622 46056
rect 31662 46044 31668 46056
rect 31720 46084 31726 46096
rect 31720 46056 45692 46084
rect 31720 46044 31726 46056
rect 1394 45948 1400 45960
rect 1355 45920 1400 45948
rect 1394 45908 1400 45920
rect 1452 45908 1458 45960
rect 2314 45948 2320 45960
rect 2275 45920 2320 45948
rect 2314 45908 2320 45920
rect 2372 45908 2378 45960
rect 3142 45948 3148 45960
rect 3103 45920 3148 45948
rect 3142 45908 3148 45920
rect 3200 45908 3206 45960
rect 42245 45951 42303 45957
rect 42245 45917 42257 45951
rect 42291 45917 42303 45951
rect 42245 45911 42303 45917
rect 1596 45852 6914 45880
rect 1596 45821 1624 45852
rect 1581 45815 1639 45821
rect 1581 45781 1593 45815
rect 1627 45781 1639 45815
rect 6886 45812 6914 45852
rect 21358 45812 21364 45824
rect 6886 45784 21364 45812
rect 1581 45775 1639 45781
rect 21358 45772 21364 45784
rect 21416 45772 21422 45824
rect 26418 45772 26424 45824
rect 26476 45812 26482 45824
rect 41969 45815 42027 45821
rect 41969 45812 41981 45815
rect 26476 45784 41981 45812
rect 26476 45772 26482 45784
rect 41969 45781 41981 45784
rect 42015 45812 42027 45815
rect 42260 45812 42288 45911
rect 44358 45908 44364 45960
rect 44416 45948 44422 45960
rect 45664 45957 45692 46056
rect 46750 46016 46756 46028
rect 45756 45988 46756 46016
rect 45005 45951 45063 45957
rect 45005 45948 45017 45951
rect 44416 45920 45017 45948
rect 44416 45908 44422 45920
rect 45005 45917 45017 45920
rect 45051 45917 45063 45951
rect 45005 45911 45063 45917
rect 45649 45951 45707 45957
rect 45649 45917 45661 45951
rect 45695 45917 45707 45951
rect 45649 45911 45707 45917
rect 45020 45880 45048 45911
rect 45756 45880 45784 45988
rect 46750 45976 46756 45988
rect 46808 45976 46814 46028
rect 48130 46016 48136 46028
rect 48091 45988 48136 46016
rect 48130 45976 48136 45988
rect 48188 45976 48194 46028
rect 46290 45948 46296 45960
rect 46251 45920 46296 45948
rect 46290 45908 46296 45920
rect 46348 45908 46354 45960
rect 45020 45852 45784 45880
rect 46477 45883 46535 45889
rect 46477 45849 46489 45883
rect 46523 45880 46535 45883
rect 47670 45880 47676 45892
rect 46523 45852 47676 45880
rect 46523 45849 46535 45852
rect 46477 45843 46535 45849
rect 47670 45840 47676 45852
rect 47728 45840 47734 45892
rect 47210 45812 47216 45824
rect 42015 45784 47216 45812
rect 42015 45781 42027 45784
rect 41969 45775 42027 45781
rect 47210 45772 47216 45784
rect 47268 45772 47274 45824
rect 1104 45722 48852 45744
rect 1104 45670 19574 45722
rect 19626 45670 19638 45722
rect 19690 45670 19702 45722
rect 19754 45670 19766 45722
rect 19818 45670 19830 45722
rect 19882 45670 48852 45722
rect 1104 45648 48852 45670
rect 3142 45540 3148 45552
rect 1780 45512 3148 45540
rect 1780 45481 1808 45512
rect 3142 45500 3148 45512
rect 3200 45500 3206 45552
rect 28258 45500 28264 45552
rect 28316 45540 28322 45552
rect 28316 45512 47624 45540
rect 28316 45500 28322 45512
rect 1765 45475 1823 45481
rect 1765 45441 1777 45475
rect 1811 45441 1823 45475
rect 1765 45435 1823 45441
rect 44085 45475 44143 45481
rect 44085 45441 44097 45475
rect 44131 45472 44143 45475
rect 44174 45472 44180 45484
rect 44131 45444 44180 45472
rect 44131 45441 44143 45444
rect 44085 45435 44143 45441
rect 44174 45432 44180 45444
rect 44232 45432 44238 45484
rect 44726 45472 44732 45484
rect 44687 45444 44732 45472
rect 44726 45432 44732 45444
rect 44784 45432 44790 45484
rect 47596 45481 47624 45512
rect 47670 45500 47676 45552
rect 47728 45540 47734 45552
rect 47728 45512 47773 45540
rect 47728 45500 47734 45512
rect 47581 45475 47639 45481
rect 47581 45441 47593 45475
rect 47627 45441 47639 45475
rect 47581 45435 47639 45441
rect 1946 45404 1952 45416
rect 1907 45376 1952 45404
rect 1946 45364 1952 45376
rect 2004 45364 2010 45416
rect 2774 45404 2780 45416
rect 2735 45376 2780 45404
rect 2774 45364 2780 45376
rect 2832 45364 2838 45416
rect 45186 45404 45192 45416
rect 45147 45376 45192 45404
rect 45186 45364 45192 45376
rect 45244 45364 45250 45416
rect 45373 45407 45431 45413
rect 45373 45373 45385 45407
rect 45419 45373 45431 45407
rect 46842 45404 46848 45416
rect 46803 45376 46848 45404
rect 45373 45367 45431 45373
rect 45388 45336 45416 45367
rect 46842 45364 46848 45376
rect 46900 45364 46906 45416
rect 47670 45336 47676 45348
rect 45388 45308 47676 45336
rect 47670 45296 47676 45308
rect 47728 45296 47734 45348
rect 1104 45178 48852 45200
rect 1104 45126 4214 45178
rect 4266 45126 4278 45178
rect 4330 45126 4342 45178
rect 4394 45126 4406 45178
rect 4458 45126 4470 45178
rect 4522 45126 34934 45178
rect 34986 45126 34998 45178
rect 35050 45126 35062 45178
rect 35114 45126 35126 45178
rect 35178 45126 35190 45178
rect 35242 45126 48852 45178
rect 1104 45104 48852 45126
rect 45186 45064 45192 45076
rect 45147 45036 45192 45064
rect 45186 45024 45192 45036
rect 45244 45024 45250 45076
rect 45554 45024 45560 45076
rect 45612 45024 45618 45076
rect 45741 45067 45799 45073
rect 45741 45033 45753 45067
rect 45787 45064 45799 45067
rect 45830 45064 45836 45076
rect 45787 45036 45836 45064
rect 45787 45033 45799 45036
rect 45741 45027 45799 45033
rect 45830 45024 45836 45036
rect 45888 45024 45894 45076
rect 2774 44928 2780 44940
rect 2735 44900 2780 44928
rect 2774 44888 2780 44900
rect 2832 44888 2838 44940
rect 1397 44863 1455 44869
rect 1397 44829 1409 44863
rect 1443 44829 1455 44863
rect 45572 44860 45600 45024
rect 46293 44931 46351 44937
rect 46293 44897 46305 44931
rect 46339 44928 46351 44931
rect 46750 44928 46756 44940
rect 46339 44900 46756 44928
rect 46339 44897 46351 44900
rect 46293 44891 46351 44897
rect 46750 44888 46756 44900
rect 46808 44888 46814 44940
rect 48130 44928 48136 44940
rect 48091 44900 48136 44928
rect 48130 44888 48136 44900
rect 48188 44888 48194 44940
rect 45649 44863 45707 44869
rect 45649 44860 45661 44863
rect 45572 44832 45661 44860
rect 1397 44823 1455 44829
rect 45649 44829 45661 44832
rect 45695 44860 45707 44863
rect 45922 44860 45928 44872
rect 45695 44832 45928 44860
rect 45695 44829 45707 44832
rect 45649 44823 45707 44829
rect 1412 44724 1440 44823
rect 45922 44820 45928 44832
rect 45980 44820 45986 44872
rect 1581 44795 1639 44801
rect 1581 44761 1593 44795
rect 1627 44792 1639 44795
rect 3418 44792 3424 44804
rect 1627 44764 3424 44792
rect 1627 44761 1639 44764
rect 1581 44755 1639 44761
rect 3418 44752 3424 44764
rect 3476 44752 3482 44804
rect 46477 44795 46535 44801
rect 46477 44761 46489 44795
rect 46523 44792 46535 44795
rect 46934 44792 46940 44804
rect 46523 44764 46940 44792
rect 46523 44761 46535 44764
rect 46477 44755 46535 44761
rect 46934 44752 46940 44764
rect 46992 44752 46998 44804
rect 2866 44724 2872 44736
rect 1412 44696 2872 44724
rect 2866 44684 2872 44696
rect 2924 44684 2930 44736
rect 1104 44634 48852 44656
rect 1104 44582 19574 44634
rect 19626 44582 19638 44634
rect 19690 44582 19702 44634
rect 19754 44582 19766 44634
rect 19818 44582 19830 44634
rect 19882 44582 48852 44634
rect 1104 44560 48852 44582
rect 1946 44480 1952 44532
rect 2004 44520 2010 44532
rect 2777 44523 2835 44529
rect 2777 44520 2789 44523
rect 2004 44492 2789 44520
rect 2004 44480 2010 44492
rect 2777 44489 2789 44492
rect 2823 44489 2835 44523
rect 3418 44520 3424 44532
rect 3379 44492 3424 44520
rect 2777 44483 2835 44489
rect 3418 44480 3424 44492
rect 3476 44480 3482 44532
rect 46934 44520 46940 44532
rect 46895 44492 46940 44520
rect 46934 44480 46940 44492
rect 46992 44480 46998 44532
rect 47670 44520 47676 44532
rect 47631 44492 47676 44520
rect 47670 44480 47676 44492
rect 47728 44480 47734 44532
rect 1854 44384 1860 44396
rect 1815 44356 1860 44384
rect 1854 44344 1860 44356
rect 1912 44344 1918 44396
rect 2222 44344 2228 44396
rect 2280 44384 2286 44396
rect 2685 44387 2743 44393
rect 2685 44384 2697 44387
rect 2280 44356 2697 44384
rect 2280 44344 2286 44356
rect 2685 44353 2697 44356
rect 2731 44353 2743 44387
rect 3326 44384 3332 44396
rect 3287 44356 3332 44384
rect 2685 44347 2743 44353
rect 3326 44344 3332 44356
rect 3384 44344 3390 44396
rect 45094 44344 45100 44396
rect 45152 44384 45158 44396
rect 45281 44387 45339 44393
rect 45281 44384 45293 44387
rect 45152 44356 45293 44384
rect 45152 44344 45158 44356
rect 45281 44353 45293 44356
rect 45327 44353 45339 44387
rect 45281 44347 45339 44353
rect 46290 44344 46296 44396
rect 46348 44384 46354 44396
rect 46385 44387 46443 44393
rect 46385 44384 46397 44387
rect 46348 44356 46397 44384
rect 46348 44344 46354 44356
rect 46385 44353 46397 44356
rect 46431 44353 46443 44387
rect 46385 44347 46443 44353
rect 46566 44344 46572 44396
rect 46624 44384 46630 44396
rect 46845 44387 46903 44393
rect 46845 44384 46857 44387
rect 46624 44356 46857 44384
rect 46624 44344 46630 44356
rect 46845 44353 46857 44356
rect 46891 44353 46903 44387
rect 46845 44347 46903 44353
rect 47486 44344 47492 44396
rect 47544 44384 47550 44396
rect 47581 44387 47639 44393
rect 47581 44384 47593 44387
rect 47544 44356 47593 44384
rect 47544 44344 47550 44356
rect 47581 44353 47593 44356
rect 47627 44353 47639 44387
rect 47581 44347 47639 44353
rect 36538 44276 36544 44328
rect 36596 44316 36602 44328
rect 45554 44316 45560 44328
rect 36596 44288 45560 44316
rect 36596 44276 36602 44288
rect 45554 44276 45560 44288
rect 45612 44276 45618 44328
rect 20346 44208 20352 44260
rect 20404 44248 20410 44260
rect 20530 44248 20536 44260
rect 20404 44220 20536 44248
rect 20404 44208 20410 44220
rect 20530 44208 20536 44220
rect 20588 44208 20594 44260
rect 43438 44208 43444 44260
rect 43496 44248 43502 44260
rect 46014 44248 46020 44260
rect 43496 44220 46020 44248
rect 43496 44208 43502 44220
rect 46014 44208 46020 44220
rect 46072 44208 46078 44260
rect 2130 44180 2136 44192
rect 2091 44152 2136 44180
rect 2130 44140 2136 44152
rect 2188 44140 2194 44192
rect 45646 44140 45652 44192
rect 45704 44180 45710 44192
rect 45922 44180 45928 44192
rect 45704 44152 45928 44180
rect 45704 44140 45710 44152
rect 45922 44140 45928 44152
rect 45980 44140 45986 44192
rect 1104 44090 48852 44112
rect 1104 44038 4214 44090
rect 4266 44038 4278 44090
rect 4330 44038 4342 44090
rect 4394 44038 4406 44090
rect 4458 44038 4470 44090
rect 4522 44038 34934 44090
rect 34986 44038 34998 44090
rect 35050 44038 35062 44090
rect 35114 44038 35126 44090
rect 35178 44038 35190 44090
rect 35242 44038 48852 44090
rect 1104 44016 48852 44038
rect 2866 43976 2872 43988
rect 2827 43948 2872 43976
rect 2866 43936 2872 43948
rect 2924 43936 2930 43988
rect 46750 43976 46756 43988
rect 46711 43948 46756 43976
rect 46750 43936 46756 43948
rect 46808 43936 46814 43988
rect 46658 43868 46664 43920
rect 46716 43908 46722 43920
rect 47397 43911 47455 43917
rect 47397 43908 47409 43911
rect 46716 43880 47409 43908
rect 46716 43868 46722 43880
rect 47397 43877 47409 43880
rect 47443 43877 47455 43911
rect 47397 43871 47455 43877
rect 21910 43800 21916 43852
rect 21968 43840 21974 43852
rect 27709 43843 27767 43849
rect 27709 43840 27721 43843
rect 21968 43812 27721 43840
rect 21968 43800 21974 43812
rect 27709 43809 27721 43812
rect 27755 43840 27767 43843
rect 27755 43812 28994 43840
rect 27755 43809 27767 43812
rect 27709 43803 27767 43809
rect 7742 43732 7748 43784
rect 7800 43772 7806 43784
rect 26694 43772 26700 43784
rect 7800 43744 26700 43772
rect 7800 43732 7806 43744
rect 26694 43732 26700 43744
rect 26752 43772 26758 43784
rect 27249 43775 27307 43781
rect 27249 43772 27261 43775
rect 26752 43744 27261 43772
rect 26752 43732 26758 43744
rect 27249 43741 27261 43744
rect 27295 43741 27307 43775
rect 27249 43735 27307 43741
rect 1854 43704 1860 43716
rect 1815 43676 1860 43704
rect 1854 43664 1860 43676
rect 1912 43664 1918 43716
rect 28966 43704 28994 43812
rect 47854 43772 47860 43784
rect 47815 43744 47860 43772
rect 47854 43732 47860 43744
rect 47912 43732 47918 43784
rect 47486 43704 47492 43716
rect 28966 43676 47492 43704
rect 47486 43664 47492 43676
rect 47544 43704 47550 43716
rect 48222 43704 48228 43716
rect 47544 43676 48228 43704
rect 47544 43664 47550 43676
rect 48222 43664 48228 43676
rect 48280 43664 48286 43716
rect 1670 43596 1676 43648
rect 1728 43636 1734 43648
rect 1949 43639 2007 43645
rect 1949 43636 1961 43639
rect 1728 43608 1961 43636
rect 1728 43596 1734 43608
rect 1949 43605 1961 43608
rect 1995 43605 2007 43639
rect 1949 43599 2007 43605
rect 46934 43596 46940 43648
rect 46992 43636 46998 43648
rect 48041 43639 48099 43645
rect 48041 43636 48053 43639
rect 46992 43608 48053 43636
rect 46992 43596 46998 43608
rect 48041 43605 48053 43608
rect 48087 43605 48099 43639
rect 48041 43599 48099 43605
rect 1104 43546 48852 43568
rect 1104 43494 19574 43546
rect 19626 43494 19638 43546
rect 19690 43494 19702 43546
rect 19754 43494 19766 43546
rect 19818 43494 19830 43546
rect 19882 43494 48852 43546
rect 1104 43472 48852 43494
rect 23382 43392 23388 43444
rect 23440 43432 23446 43444
rect 47302 43432 47308 43444
rect 23440 43404 47308 43432
rect 23440 43392 23446 43404
rect 47302 43392 47308 43404
rect 47360 43392 47366 43444
rect 47946 43296 47952 43308
rect 47907 43268 47952 43296
rect 47946 43256 47952 43268
rect 48004 43256 48010 43308
rect 47026 43092 47032 43104
rect 46987 43064 47032 43092
rect 47026 43052 47032 43064
rect 47084 43052 47090 43104
rect 48038 43092 48044 43104
rect 47999 43064 48044 43092
rect 48038 43052 48044 43064
rect 48096 43052 48102 43104
rect 1104 43002 48852 43024
rect 1104 42950 4214 43002
rect 4266 42950 4278 43002
rect 4330 42950 4342 43002
rect 4394 42950 4406 43002
rect 4458 42950 4470 43002
rect 4522 42950 34934 43002
rect 34986 42950 34998 43002
rect 35050 42950 35062 43002
rect 35114 42950 35126 43002
rect 35178 42950 35190 43002
rect 35242 42950 48852 43002
rect 1104 42928 48852 42950
rect 46293 42755 46351 42761
rect 46293 42721 46305 42755
rect 46339 42752 46351 42755
rect 47026 42752 47032 42764
rect 46339 42724 47032 42752
rect 46339 42721 46351 42724
rect 46293 42715 46351 42721
rect 47026 42712 47032 42724
rect 47084 42712 47090 42764
rect 48130 42752 48136 42764
rect 48091 42724 48136 42752
rect 48130 42712 48136 42724
rect 48188 42712 48194 42764
rect 46474 42616 46480 42628
rect 46435 42588 46480 42616
rect 46474 42576 46480 42588
rect 46532 42576 46538 42628
rect 1104 42458 48852 42480
rect 1104 42406 19574 42458
rect 19626 42406 19638 42458
rect 19690 42406 19702 42458
rect 19754 42406 19766 42458
rect 19818 42406 19830 42458
rect 19882 42406 48852 42458
rect 1104 42384 48852 42406
rect 45738 42236 45744 42288
rect 45796 42276 45802 42288
rect 46474 42276 46480 42288
rect 45796 42248 46480 42276
rect 45796 42236 45802 42248
rect 46474 42236 46480 42248
rect 46532 42276 46538 42288
rect 47581 42279 47639 42285
rect 47581 42276 47593 42279
rect 46532 42248 47593 42276
rect 46532 42236 46538 42248
rect 47581 42245 47593 42248
rect 47627 42245 47639 42279
rect 47581 42239 47639 42245
rect 22741 42211 22799 42217
rect 22741 42177 22753 42211
rect 22787 42177 22799 42211
rect 22922 42208 22928 42220
rect 22883 42180 22928 42208
rect 22741 42171 22799 42177
rect 20714 42100 20720 42152
rect 20772 42140 20778 42152
rect 22756 42140 22784 42171
rect 22922 42168 22928 42180
rect 22980 42168 22986 42220
rect 23017 42211 23075 42217
rect 23017 42177 23029 42211
rect 23063 42208 23075 42211
rect 24578 42208 24584 42220
rect 23063 42180 24584 42208
rect 23063 42177 23075 42180
rect 23017 42171 23075 42177
rect 24578 42168 24584 42180
rect 24636 42168 24642 42220
rect 47210 42168 47216 42220
rect 47268 42208 47274 42220
rect 47854 42208 47860 42220
rect 47268 42180 47860 42208
rect 47268 42168 47274 42180
rect 47854 42168 47860 42180
rect 47912 42168 47918 42220
rect 25866 42140 25872 42152
rect 20772 42112 25872 42140
rect 20772 42100 20778 42112
rect 25866 42100 25872 42112
rect 25924 42100 25930 42152
rect 1394 41964 1400 42016
rect 1452 42004 1458 42016
rect 2041 42007 2099 42013
rect 2041 42004 2053 42007
rect 1452 41976 2053 42004
rect 1452 41964 1458 41976
rect 2041 41973 2053 41976
rect 2087 41973 2099 42007
rect 2041 41967 2099 41973
rect 22557 42007 22615 42013
rect 22557 41973 22569 42007
rect 22603 42004 22615 42007
rect 23566 42004 23572 42016
rect 22603 41976 23572 42004
rect 22603 41973 22615 41976
rect 22557 41967 22615 41973
rect 23566 41964 23572 41976
rect 23624 41964 23630 42016
rect 1104 41914 48852 41936
rect 1104 41862 4214 41914
rect 4266 41862 4278 41914
rect 4330 41862 4342 41914
rect 4394 41862 4406 41914
rect 4458 41862 4470 41914
rect 4522 41862 34934 41914
rect 34986 41862 34998 41914
rect 35050 41862 35062 41914
rect 35114 41862 35126 41914
rect 35178 41862 35190 41914
rect 35242 41862 48852 41914
rect 1104 41840 48852 41862
rect 48038 41732 48044 41744
rect 23400 41704 48044 41732
rect 1394 41664 1400 41676
rect 1355 41636 1400 41664
rect 1394 41624 1400 41636
rect 1452 41624 1458 41676
rect 1854 41664 1860 41676
rect 1815 41636 1860 41664
rect 1854 41624 1860 41636
rect 1912 41624 1918 41676
rect 19245 41599 19303 41605
rect 19245 41565 19257 41599
rect 19291 41596 19303 41599
rect 19334 41596 19340 41608
rect 19291 41568 19340 41596
rect 19291 41565 19303 41568
rect 19245 41559 19303 41565
rect 19334 41556 19340 41568
rect 19392 41596 19398 41608
rect 23400 41605 23428 41704
rect 48038 41692 48044 41704
rect 48096 41692 48102 41744
rect 46293 41667 46351 41673
rect 46293 41633 46305 41667
rect 46339 41664 46351 41667
rect 47670 41664 47676 41676
rect 46339 41636 47676 41664
rect 46339 41633 46351 41636
rect 46293 41627 46351 41633
rect 47670 41624 47676 41636
rect 47728 41624 47734 41676
rect 21269 41599 21327 41605
rect 21269 41596 21281 41599
rect 19392 41568 21281 41596
rect 19392 41556 19398 41568
rect 21269 41565 21281 41568
rect 21315 41565 21327 41599
rect 21269 41559 21327 41565
rect 23385 41599 23443 41605
rect 23385 41565 23397 41599
rect 23431 41565 23443 41599
rect 23385 41559 23443 41565
rect 23477 41599 23535 41605
rect 23477 41565 23489 41599
rect 23523 41565 23535 41599
rect 23477 41559 23535 41565
rect 1578 41528 1584 41540
rect 1539 41500 1584 41528
rect 1578 41488 1584 41500
rect 1636 41488 1642 41540
rect 19512 41531 19570 41537
rect 19512 41497 19524 41531
rect 19558 41497 19570 41531
rect 19512 41491 19570 41497
rect 21536 41531 21594 41537
rect 21536 41497 21548 41531
rect 21582 41528 21594 41531
rect 21818 41528 21824 41540
rect 21582 41500 21824 41528
rect 21582 41497 21594 41500
rect 21536 41491 21594 41497
rect 19426 41420 19432 41472
rect 19484 41460 19490 41472
rect 19536 41460 19564 41491
rect 21818 41488 21824 41500
rect 21876 41488 21882 41540
rect 22370 41488 22376 41540
rect 22428 41528 22434 41540
rect 23014 41528 23020 41540
rect 22428 41500 23020 41528
rect 22428 41488 22434 41500
rect 23014 41488 23020 41500
rect 23072 41528 23078 41540
rect 23492 41528 23520 41559
rect 23566 41556 23572 41608
rect 23624 41596 23630 41608
rect 23750 41596 23756 41608
rect 23624 41568 23669 41596
rect 23711 41568 23756 41596
rect 23624 41556 23630 41568
rect 23750 41556 23756 41568
rect 23808 41556 23814 41608
rect 46474 41528 46480 41540
rect 23072 41500 23520 41528
rect 46435 41500 46480 41528
rect 23072 41488 23078 41500
rect 46474 41488 46480 41500
rect 46532 41488 46538 41540
rect 48130 41528 48136 41540
rect 48091 41500 48136 41528
rect 48130 41488 48136 41500
rect 48188 41488 48194 41540
rect 19484 41432 19564 41460
rect 20625 41463 20683 41469
rect 19484 41420 19490 41432
rect 20625 41429 20637 41463
rect 20671 41460 20683 41463
rect 20898 41460 20904 41472
rect 20671 41432 20904 41460
rect 20671 41429 20683 41432
rect 20625 41423 20683 41429
rect 20898 41420 20904 41432
rect 20956 41420 20962 41472
rect 22186 41420 22192 41472
rect 22244 41460 22250 41472
rect 22649 41463 22707 41469
rect 22649 41460 22661 41463
rect 22244 41432 22661 41460
rect 22244 41420 22250 41432
rect 22649 41429 22661 41432
rect 22695 41429 22707 41463
rect 22649 41423 22707 41429
rect 23109 41463 23167 41469
rect 23109 41429 23121 41463
rect 23155 41460 23167 41463
rect 23474 41460 23480 41472
rect 23155 41432 23480 41460
rect 23155 41429 23167 41432
rect 23109 41423 23167 41429
rect 23474 41420 23480 41432
rect 23532 41420 23538 41472
rect 1104 41370 48852 41392
rect 1104 41318 19574 41370
rect 19626 41318 19638 41370
rect 19690 41318 19702 41370
rect 19754 41318 19766 41370
rect 19818 41318 19830 41370
rect 19882 41318 48852 41370
rect 1104 41296 48852 41318
rect 1578 41216 1584 41268
rect 1636 41256 1642 41268
rect 2593 41259 2651 41265
rect 2593 41256 2605 41259
rect 1636 41228 2605 41256
rect 1636 41216 1642 41228
rect 2593 41225 2605 41228
rect 2639 41225 2651 41259
rect 2593 41219 2651 41225
rect 18877 41259 18935 41265
rect 18877 41225 18889 41259
rect 18923 41256 18935 41259
rect 19426 41256 19432 41268
rect 18923 41228 19432 41256
rect 18923 41225 18935 41228
rect 18877 41219 18935 41225
rect 19426 41216 19432 41228
rect 19484 41216 19490 41268
rect 21818 41256 21824 41268
rect 21779 41228 21824 41256
rect 21818 41216 21824 41228
rect 21876 41216 21882 41268
rect 22278 41256 22284 41268
rect 22112 41228 22284 41256
rect 21910 41188 21916 41200
rect 2746 41160 21916 41188
rect 1854 41120 1860 41132
rect 1815 41092 1860 41120
rect 1854 41080 1860 41092
rect 1912 41080 1918 41132
rect 2314 41080 2320 41132
rect 2372 41120 2378 41132
rect 2501 41123 2559 41129
rect 2501 41120 2513 41123
rect 2372 41092 2513 41120
rect 2372 41080 2378 41092
rect 2501 41089 2513 41092
rect 2547 41120 2559 41123
rect 2746 41120 2774 41160
rect 21910 41148 21916 41160
rect 21968 41148 21974 41200
rect 2547 41092 2774 41120
rect 2547 41089 2559 41092
rect 2501 41083 2559 41089
rect 2958 41080 2964 41132
rect 3016 41120 3022 41132
rect 19153 41123 19211 41129
rect 19153 41120 19165 41123
rect 3016 41092 19165 41120
rect 3016 41080 3022 41092
rect 19153 41089 19165 41092
rect 19199 41089 19211 41123
rect 19153 41083 19211 41089
rect 19245 41123 19303 41129
rect 19245 41089 19257 41123
rect 19291 41089 19303 41123
rect 19245 41083 19303 41089
rect 19337 41123 19395 41129
rect 19337 41089 19349 41123
rect 19383 41089 19395 41123
rect 19337 41083 19395 41089
rect 19521 41123 19579 41129
rect 19521 41089 19533 41123
rect 19567 41120 19579 41123
rect 20070 41120 20076 41132
rect 19567 41092 20076 41120
rect 19567 41089 19579 41092
rect 19521 41083 19579 41089
rect 18782 41012 18788 41064
rect 18840 41052 18846 41064
rect 19260 41052 19288 41083
rect 18840 41024 19288 41052
rect 19352 41052 19380 41083
rect 20070 41080 20076 41092
rect 20128 41080 20134 41132
rect 20165 41123 20223 41129
rect 20165 41089 20177 41123
rect 20211 41120 20223 41123
rect 20349 41123 20407 41129
rect 20211 41092 20300 41120
rect 20211 41089 20223 41092
rect 20165 41083 20223 41089
rect 19981 41055 20039 41061
rect 19981 41052 19993 41055
rect 19352 41024 19993 41052
rect 18840 41012 18846 41024
rect 19981 41021 19993 41024
rect 20027 41021 20039 41055
rect 19981 41015 20039 41021
rect 2041 40987 2099 40993
rect 2041 40953 2053 40987
rect 2087 40984 2099 40987
rect 2406 40984 2412 40996
rect 2087 40956 2412 40984
rect 2087 40953 2099 40956
rect 2041 40947 2099 40953
rect 2406 40944 2412 40956
rect 2464 40944 2470 40996
rect 20272 40984 20300 41092
rect 20349 41089 20361 41123
rect 20395 41089 20407 41123
rect 20349 41083 20407 41089
rect 20441 41123 20499 41129
rect 20441 41089 20453 41123
rect 20487 41120 20499 41123
rect 20898 41120 20904 41132
rect 20487 41092 20904 41120
rect 20487 41089 20499 41092
rect 20441 41083 20499 41089
rect 20364 41052 20392 41083
rect 20898 41080 20904 41092
rect 20956 41080 20962 41132
rect 22112 41129 22140 41228
rect 22278 41216 22284 41228
rect 22336 41216 22342 41268
rect 46474 41216 46480 41268
rect 46532 41256 46538 41268
rect 46753 41259 46811 41265
rect 46753 41256 46765 41259
rect 46532 41228 46765 41256
rect 46532 41216 46538 41228
rect 46753 41225 46765 41228
rect 46799 41225 46811 41259
rect 46753 41219 46811 41225
rect 23474 41197 23480 41200
rect 23468 41188 23480 41197
rect 23435 41160 23480 41188
rect 23468 41151 23480 41160
rect 23474 41148 23480 41151
rect 23532 41148 23538 41200
rect 22097 41123 22155 41129
rect 22097 41089 22109 41123
rect 22143 41089 22155 41123
rect 22097 41083 22155 41089
rect 22189 41123 22247 41129
rect 22189 41089 22201 41123
rect 22235 41089 22247 41123
rect 22189 41083 22247 41089
rect 20806 41052 20812 41064
rect 20364 41024 20812 41052
rect 20806 41012 20812 41024
rect 20864 41012 20870 41064
rect 22204 41052 22232 41083
rect 22278 41080 22284 41132
rect 22336 41120 22342 41132
rect 22465 41123 22523 41129
rect 22336 41092 22381 41120
rect 22336 41080 22342 41092
rect 22465 41089 22477 41123
rect 22511 41120 22523 41123
rect 23750 41120 23756 41132
rect 22511 41092 23756 41120
rect 22511 41089 22523 41092
rect 22465 41083 22523 41089
rect 23750 41080 23756 41092
rect 23808 41080 23814 41132
rect 46658 41120 46664 41132
rect 46619 41092 46664 41120
rect 46658 41080 46664 41092
rect 46716 41080 46722 41132
rect 47670 41080 47676 41132
rect 47728 41120 47734 41132
rect 47765 41123 47823 41129
rect 47765 41120 47777 41123
rect 47728 41092 47777 41120
rect 47728 41080 47734 41092
rect 47765 41089 47777 41092
rect 47811 41089 47823 41123
rect 47765 41083 47823 41089
rect 22370 41052 22376 41064
rect 22204 41024 22376 41052
rect 22370 41012 22376 41024
rect 22428 41012 22434 41064
rect 23198 41052 23204 41064
rect 23159 41024 23204 41052
rect 23198 41012 23204 41024
rect 23256 41012 23262 41064
rect 20714 40984 20720 40996
rect 20272 40956 20720 40984
rect 19978 40876 19984 40928
rect 20036 40916 20042 40928
rect 20272 40916 20300 40956
rect 20714 40944 20720 40956
rect 20772 40944 20778 40996
rect 20036 40888 20300 40916
rect 24581 40919 24639 40925
rect 20036 40876 20042 40888
rect 24581 40885 24593 40919
rect 24627 40916 24639 40919
rect 24670 40916 24676 40928
rect 24627 40888 24676 40916
rect 24627 40885 24639 40888
rect 24581 40879 24639 40885
rect 24670 40876 24676 40888
rect 24728 40876 24734 40928
rect 1104 40826 48852 40848
rect 1104 40774 4214 40826
rect 4266 40774 4278 40826
rect 4330 40774 4342 40826
rect 4394 40774 4406 40826
rect 4458 40774 4470 40826
rect 4522 40774 34934 40826
rect 34986 40774 34998 40826
rect 35050 40774 35062 40826
rect 35114 40774 35126 40826
rect 35178 40774 35190 40826
rect 35242 40774 48852 40826
rect 1104 40752 48852 40774
rect 21637 40715 21695 40721
rect 21637 40681 21649 40715
rect 21683 40712 21695 40715
rect 22278 40712 22284 40724
rect 21683 40684 22284 40712
rect 21683 40681 21695 40684
rect 21637 40675 21695 40681
rect 22278 40672 22284 40684
rect 22336 40672 22342 40724
rect 29822 40712 29828 40724
rect 22572 40684 29828 40712
rect 19628 40548 21864 40576
rect 1394 40508 1400 40520
rect 1355 40480 1400 40508
rect 1394 40468 1400 40480
rect 1452 40468 1458 40520
rect 18598 40468 18604 40520
rect 18656 40508 18662 40520
rect 19628 40517 19656 40548
rect 19613 40511 19671 40517
rect 19613 40508 19625 40511
rect 18656 40480 19625 40508
rect 18656 40468 18662 40480
rect 19613 40477 19625 40480
rect 19659 40477 19671 40511
rect 19613 40471 19671 40477
rect 19889 40511 19947 40517
rect 19889 40477 19901 40511
rect 19935 40508 19947 40511
rect 20438 40508 20444 40520
rect 19935 40480 20444 40508
rect 19935 40477 19947 40480
rect 19889 40471 19947 40477
rect 20438 40468 20444 40480
rect 20496 40468 20502 40520
rect 21836 40517 21864 40548
rect 21821 40511 21879 40517
rect 21821 40477 21833 40511
rect 21867 40477 21879 40511
rect 21821 40471 21879 40477
rect 21836 40440 21864 40471
rect 22094 40468 22100 40520
rect 22152 40508 22158 40520
rect 22572 40508 22600 40684
rect 29822 40672 29828 40684
rect 29880 40672 29886 40724
rect 22646 40536 22652 40588
rect 22704 40576 22710 40588
rect 23198 40576 23204 40588
rect 22704 40548 23204 40576
rect 22704 40536 22710 40548
rect 23198 40536 23204 40548
rect 23256 40576 23262 40588
rect 24489 40579 24547 40585
rect 24489 40576 24501 40579
rect 23256 40548 24501 40576
rect 23256 40536 23262 40548
rect 24489 40545 24501 40548
rect 24535 40545 24547 40579
rect 47302 40576 47308 40588
rect 47263 40548 47308 40576
rect 24489 40539 24547 40545
rect 47302 40536 47308 40548
rect 47360 40536 47366 40588
rect 22741 40511 22799 40517
rect 22741 40508 22753 40511
rect 22152 40480 22197 40508
rect 22480 40480 22753 40508
rect 22152 40468 22158 40480
rect 22480 40440 22508 40480
rect 22741 40477 22753 40480
rect 22787 40477 22799 40511
rect 22922 40508 22928 40520
rect 22883 40480 22928 40508
rect 22741 40471 22799 40477
rect 22922 40468 22928 40480
rect 22980 40468 22986 40520
rect 23017 40511 23075 40517
rect 23017 40477 23029 40511
rect 23063 40508 23075 40511
rect 23063 40480 24900 40508
rect 23063 40477 23075 40480
rect 23017 40471 23075 40477
rect 24872 40452 24900 40480
rect 47394 40468 47400 40520
rect 47452 40508 47458 40520
rect 47581 40511 47639 40517
rect 47581 40508 47593 40511
rect 47452 40480 47593 40508
rect 47452 40468 47458 40480
rect 47581 40477 47593 40480
rect 47627 40477 47639 40511
rect 47581 40471 47639 40477
rect 21836 40412 22508 40440
rect 22557 40443 22615 40449
rect 22557 40409 22569 40443
rect 22603 40440 22615 40443
rect 23106 40440 23112 40452
rect 22603 40412 23112 40440
rect 22603 40409 22615 40412
rect 22557 40403 22615 40409
rect 23106 40400 23112 40412
rect 23164 40400 23170 40452
rect 24578 40400 24584 40452
rect 24636 40440 24642 40452
rect 24734 40443 24792 40449
rect 24734 40440 24746 40443
rect 24636 40412 24746 40440
rect 24636 40400 24642 40412
rect 24734 40409 24746 40412
rect 24780 40409 24792 40443
rect 24734 40403 24792 40409
rect 24854 40400 24860 40452
rect 24912 40400 24918 40452
rect 1578 40372 1584 40384
rect 1539 40344 1584 40372
rect 1578 40332 1584 40344
rect 1636 40332 1642 40384
rect 19426 40372 19432 40384
rect 19387 40344 19432 40372
rect 19426 40332 19432 40344
rect 19484 40332 19490 40384
rect 19797 40375 19855 40381
rect 19797 40341 19809 40375
rect 19843 40372 19855 40375
rect 20806 40372 20812 40384
rect 19843 40344 20812 40372
rect 19843 40341 19855 40344
rect 19797 40335 19855 40341
rect 20806 40332 20812 40344
rect 20864 40372 20870 40384
rect 22005 40375 22063 40381
rect 22005 40372 22017 40375
rect 20864 40344 22017 40372
rect 20864 40332 20870 40344
rect 22005 40341 22017 40344
rect 22051 40372 22063 40375
rect 22922 40372 22928 40384
rect 22051 40344 22928 40372
rect 22051 40341 22063 40344
rect 22005 40335 22063 40341
rect 22922 40332 22928 40344
rect 22980 40332 22986 40384
rect 24486 40332 24492 40384
rect 24544 40372 24550 40384
rect 25869 40375 25927 40381
rect 25869 40372 25881 40375
rect 24544 40344 25881 40372
rect 24544 40332 24550 40344
rect 25869 40341 25881 40344
rect 25915 40341 25927 40375
rect 25869 40335 25927 40341
rect 1104 40282 48852 40304
rect 1104 40230 19574 40282
rect 19626 40230 19638 40282
rect 19690 40230 19702 40282
rect 19754 40230 19766 40282
rect 19818 40230 19830 40282
rect 19882 40230 48852 40282
rect 1104 40208 48852 40230
rect 20438 40168 20444 40180
rect 20351 40140 20444 40168
rect 20438 40128 20444 40140
rect 20496 40168 20502 40180
rect 22922 40168 22928 40180
rect 20496 40140 22928 40168
rect 20496 40128 20502 40140
rect 22922 40128 22928 40140
rect 22980 40128 22986 40180
rect 24578 40168 24584 40180
rect 24539 40140 24584 40168
rect 24578 40128 24584 40140
rect 24636 40128 24642 40180
rect 26053 40171 26111 40177
rect 26053 40137 26065 40171
rect 26099 40168 26111 40171
rect 26602 40168 26608 40180
rect 26099 40140 26608 40168
rect 26099 40137 26111 40140
rect 26053 40131 26111 40137
rect 26602 40128 26608 40140
rect 26660 40128 26666 40180
rect 26973 40171 27031 40177
rect 26973 40137 26985 40171
rect 27019 40168 27031 40171
rect 27019 40140 28212 40168
rect 27019 40137 27031 40140
rect 26973 40131 27031 40137
rect 19886 40060 19892 40112
rect 19944 40100 19950 40112
rect 20070 40100 20076 40112
rect 19944 40072 20076 40100
rect 19944 40060 19950 40072
rect 20070 40060 20076 40072
rect 20128 40100 20134 40112
rect 23750 40100 23756 40112
rect 20128 40072 23756 40100
rect 20128 40060 20134 40072
rect 23750 40060 23756 40072
rect 23808 40060 23814 40112
rect 25314 40100 25320 40112
rect 24964 40072 25320 40100
rect 18417 40035 18475 40041
rect 18417 40001 18429 40035
rect 18463 40032 18475 40035
rect 18506 40032 18512 40044
rect 18463 40004 18512 40032
rect 18463 40001 18475 40004
rect 18417 39995 18475 40001
rect 18506 39992 18512 40004
rect 18564 39992 18570 40044
rect 19150 39992 19156 40044
rect 19208 40032 19214 40044
rect 19317 40035 19375 40041
rect 19317 40032 19329 40035
rect 19208 40004 19329 40032
rect 19208 39992 19214 40004
rect 19317 40001 19329 40004
rect 19363 40001 19375 40035
rect 19317 39995 19375 40001
rect 22830 39992 22836 40044
rect 22888 40032 22894 40044
rect 22997 40035 23055 40041
rect 22997 40032 23009 40035
rect 22888 40004 23009 40032
rect 22888 39992 22894 40004
rect 22997 40001 23009 40004
rect 23043 40001 23055 40035
rect 22997 39995 23055 40001
rect 24118 39992 24124 40044
rect 24176 40032 24182 40044
rect 24964 40041 24992 40072
rect 25314 40060 25320 40072
rect 25372 40060 25378 40112
rect 27338 40100 27344 40112
rect 25700 40072 26280 40100
rect 27299 40072 27344 40100
rect 24857 40035 24915 40041
rect 24857 40032 24869 40035
rect 24176 40004 24869 40032
rect 24176 39992 24182 40004
rect 24857 40001 24869 40004
rect 24903 40001 24915 40035
rect 24857 39995 24915 40001
rect 24949 40035 25007 40041
rect 24949 40001 24961 40035
rect 24995 40001 25007 40035
rect 24949 39995 25007 40001
rect 25038 39992 25044 40044
rect 25096 40032 25102 40044
rect 25225 40035 25283 40041
rect 25096 40004 25141 40032
rect 25096 39992 25102 40004
rect 25225 40001 25237 40035
rect 25271 40032 25283 40035
rect 25700 40032 25728 40072
rect 25866 40032 25872 40044
rect 25271 40004 25728 40032
rect 25827 40004 25872 40032
rect 25271 40001 25283 40004
rect 25225 39995 25283 40001
rect 19061 39967 19119 39973
rect 19061 39933 19073 39967
rect 19107 39933 19119 39967
rect 19061 39927 19119 39933
rect 18601 39899 18659 39905
rect 18601 39865 18613 39899
rect 18647 39896 18659 39899
rect 18782 39896 18788 39908
rect 18647 39868 18788 39896
rect 18647 39865 18659 39868
rect 18601 39859 18659 39865
rect 18782 39856 18788 39868
rect 18840 39856 18846 39908
rect 19076 39828 19104 39927
rect 22186 39924 22192 39976
rect 22244 39964 22250 39976
rect 22646 39964 22652 39976
rect 22244 39936 22652 39964
rect 22244 39924 22250 39936
rect 22646 39924 22652 39936
rect 22704 39964 22710 39976
rect 22741 39967 22799 39973
rect 22741 39964 22753 39967
rect 22704 39936 22753 39964
rect 22704 39924 22710 39936
rect 22741 39933 22753 39936
rect 22787 39933 22799 39967
rect 22741 39927 22799 39933
rect 23842 39924 23848 39976
rect 23900 39964 23906 39976
rect 25240 39964 25268 39995
rect 25866 39992 25872 40004
rect 25924 39992 25930 40044
rect 26145 40035 26203 40041
rect 26145 40001 26157 40035
rect 26191 40001 26203 40035
rect 26252 40032 26280 40072
rect 27338 40060 27344 40072
rect 27396 40060 27402 40112
rect 28184 40109 28212 40140
rect 28169 40103 28227 40109
rect 28169 40069 28181 40103
rect 28215 40069 28227 40103
rect 28169 40063 28227 40069
rect 28353 40103 28411 40109
rect 28353 40069 28365 40103
rect 28399 40069 28411 40103
rect 28353 40063 28411 40069
rect 26252 40004 27752 40032
rect 26145 39995 26203 40001
rect 23900 39936 25268 39964
rect 23900 39924 23906 39936
rect 25774 39924 25780 39976
rect 25832 39964 25838 39976
rect 26160 39964 26188 39995
rect 25832 39936 26188 39964
rect 27433 39967 27491 39973
rect 25832 39924 25838 39936
rect 27433 39933 27445 39967
rect 27479 39933 27491 39967
rect 27433 39927 27491 39933
rect 20622 39896 20628 39908
rect 19996 39868 20628 39896
rect 19334 39828 19340 39840
rect 19076 39800 19340 39828
rect 19334 39788 19340 39800
rect 19392 39828 19398 39840
rect 19996 39828 20024 39868
rect 20622 39856 20628 39868
rect 20680 39856 20686 39908
rect 24946 39856 24952 39908
rect 25004 39896 25010 39908
rect 27448 39896 27476 39927
rect 27522 39924 27528 39976
rect 27580 39964 27586 39976
rect 27724 39964 27752 40004
rect 28074 39992 28080 40044
rect 28132 40032 28138 40044
rect 28368 40032 28396 40063
rect 28132 40004 28396 40032
rect 28132 39992 28138 40004
rect 43622 39992 43628 40044
rect 43680 40032 43686 40044
rect 47486 40032 47492 40044
rect 43680 40004 47492 40032
rect 43680 39992 43686 40004
rect 47486 39992 47492 40004
rect 47544 40032 47550 40044
rect 47581 40035 47639 40041
rect 47581 40032 47593 40035
rect 47544 40004 47593 40032
rect 47544 39992 47550 40004
rect 47581 40001 47593 40004
rect 47627 40001 47639 40035
rect 47581 39995 47639 40001
rect 28994 39964 29000 39976
rect 27580 39936 27625 39964
rect 27724 39936 29000 39964
rect 27580 39924 27586 39936
rect 28994 39924 29000 39936
rect 29052 39924 29058 39976
rect 25004 39868 27476 39896
rect 25004 39856 25010 39868
rect 19392 39800 20024 39828
rect 24121 39831 24179 39837
rect 19392 39788 19398 39800
rect 24121 39797 24133 39831
rect 24167 39828 24179 39831
rect 24854 39828 24860 39840
rect 24167 39800 24860 39828
rect 24167 39797 24179 39800
rect 24121 39791 24179 39797
rect 24854 39788 24860 39800
rect 24912 39788 24918 39840
rect 25685 39831 25743 39837
rect 25685 39797 25697 39831
rect 25731 39828 25743 39831
rect 26142 39828 26148 39840
rect 25731 39800 26148 39828
rect 25731 39797 25743 39800
rect 25685 39791 25743 39797
rect 26142 39788 26148 39800
rect 26200 39788 26206 39840
rect 28537 39831 28595 39837
rect 28537 39797 28549 39831
rect 28583 39828 28595 39831
rect 28902 39828 28908 39840
rect 28583 39800 28908 39828
rect 28583 39797 28595 39800
rect 28537 39791 28595 39797
rect 28902 39788 28908 39800
rect 28960 39788 28966 39840
rect 46290 39788 46296 39840
rect 46348 39828 46354 39840
rect 47029 39831 47087 39837
rect 47029 39828 47041 39831
rect 46348 39800 47041 39828
rect 46348 39788 46354 39800
rect 47029 39797 47041 39800
rect 47075 39797 47087 39831
rect 47670 39828 47676 39840
rect 47631 39800 47676 39828
rect 47029 39791 47087 39797
rect 47670 39788 47676 39800
rect 47728 39788 47734 39840
rect 1104 39738 48852 39760
rect 1104 39686 4214 39738
rect 4266 39686 4278 39738
rect 4330 39686 4342 39738
rect 4394 39686 4406 39738
rect 4458 39686 4470 39738
rect 4522 39686 34934 39738
rect 34986 39686 34998 39738
rect 35050 39686 35062 39738
rect 35114 39686 35126 39738
rect 35178 39686 35190 39738
rect 35242 39686 48852 39738
rect 1104 39664 48852 39686
rect 19150 39584 19156 39636
rect 19208 39624 19214 39636
rect 19245 39627 19303 39633
rect 19245 39624 19257 39627
rect 19208 39596 19257 39624
rect 19208 39584 19214 39596
rect 19245 39593 19257 39596
rect 19291 39593 19303 39627
rect 19245 39587 19303 39593
rect 22649 39627 22707 39633
rect 22649 39593 22661 39627
rect 22695 39624 22707 39627
rect 22830 39624 22836 39636
rect 22695 39596 22836 39624
rect 22695 39593 22707 39596
rect 22649 39587 22707 39593
rect 22830 39584 22836 39596
rect 22888 39584 22894 39636
rect 48038 39624 48044 39636
rect 24964 39596 48044 39624
rect 19426 39448 19432 39500
rect 19484 39488 19490 39500
rect 20806 39488 20812 39500
rect 19484 39460 19748 39488
rect 20767 39460 20812 39488
rect 19484 39448 19490 39460
rect 17313 39423 17371 39429
rect 17313 39389 17325 39423
rect 17359 39420 17371 39423
rect 19334 39420 19340 39432
rect 17359 39392 19340 39420
rect 17359 39389 17371 39392
rect 17313 39383 17371 39389
rect 19334 39380 19340 39392
rect 19392 39380 19398 39432
rect 19720 39429 19748 39460
rect 20806 39448 20812 39460
rect 20864 39448 20870 39500
rect 24964 39488 24992 39596
rect 48038 39584 48044 39596
rect 48096 39584 48102 39636
rect 28074 39516 28080 39568
rect 28132 39556 28138 39568
rect 28132 39528 29224 39556
rect 28132 39516 28138 39528
rect 22940 39460 24992 39488
rect 25041 39491 25099 39497
rect 19521 39423 19579 39429
rect 19521 39389 19533 39423
rect 19567 39389 19579 39423
rect 19521 39383 19579 39389
rect 19613 39423 19671 39429
rect 19613 39389 19625 39423
rect 19659 39389 19671 39423
rect 19613 39383 19671 39389
rect 19705 39423 19763 39429
rect 19705 39389 19717 39423
rect 19751 39389 19763 39423
rect 19886 39420 19892 39432
rect 19847 39392 19892 39420
rect 19705 39383 19763 39389
rect 17402 39312 17408 39364
rect 17460 39352 17466 39364
rect 17558 39355 17616 39361
rect 17558 39352 17570 39355
rect 17460 39324 17570 39352
rect 17460 39312 17466 39324
rect 17558 39321 17570 39324
rect 17604 39321 17616 39355
rect 19536 39352 19564 39383
rect 17558 39315 17616 39321
rect 18524 39324 19564 39352
rect 17218 39244 17224 39296
rect 17276 39284 17282 39296
rect 18524 39284 18552 39324
rect 18690 39284 18696 39296
rect 17276 39256 18552 39284
rect 18651 39256 18696 39284
rect 17276 39244 17282 39256
rect 18690 39244 18696 39256
rect 18748 39244 18754 39296
rect 18782 39244 18788 39296
rect 18840 39284 18846 39296
rect 19628 39284 19656 39383
rect 19886 39380 19892 39392
rect 19944 39420 19950 39432
rect 20070 39420 20076 39432
rect 19944 39392 20076 39420
rect 19944 39380 19950 39392
rect 20070 39380 20076 39392
rect 20128 39380 20134 39432
rect 20533 39423 20591 39429
rect 20533 39389 20545 39423
rect 20579 39420 20591 39423
rect 20714 39420 20720 39432
rect 20579 39392 20720 39420
rect 20579 39389 20591 39392
rect 20533 39383 20591 39389
rect 20714 39380 20720 39392
rect 20772 39380 20778 39432
rect 22940 39429 22968 39460
rect 25041 39457 25053 39491
rect 25087 39488 25099 39491
rect 26050 39488 26056 39500
rect 25087 39460 26056 39488
rect 25087 39457 25099 39460
rect 25041 39451 25099 39457
rect 26050 39448 26056 39460
rect 26108 39448 26114 39500
rect 28442 39448 28448 39500
rect 28500 39488 28506 39500
rect 28500 39460 28764 39488
rect 28500 39448 28506 39460
rect 22925 39423 22983 39429
rect 22925 39389 22937 39423
rect 22971 39389 22983 39423
rect 22925 39383 22983 39389
rect 23017 39423 23075 39429
rect 23017 39389 23029 39423
rect 23063 39389 23075 39423
rect 23017 39383 23075 39389
rect 23032 39296 23060 39383
rect 23106 39380 23112 39432
rect 23164 39420 23170 39432
rect 23293 39423 23351 39429
rect 23164 39392 23209 39420
rect 23164 39380 23170 39392
rect 23293 39389 23305 39423
rect 23339 39420 23351 39423
rect 23842 39420 23848 39432
rect 23339 39392 23848 39420
rect 23339 39389 23351 39392
rect 23293 39383 23351 39389
rect 23842 39380 23848 39392
rect 23900 39380 23906 39432
rect 24486 39380 24492 39432
rect 24544 39420 24550 39432
rect 24765 39423 24823 39429
rect 24765 39420 24777 39423
rect 24544 39392 24777 39420
rect 24544 39380 24550 39392
rect 24765 39389 24777 39392
rect 24811 39389 24823 39423
rect 24765 39383 24823 39389
rect 26237 39423 26295 39429
rect 26237 39389 26249 39423
rect 26283 39420 26295 39423
rect 28534 39420 28540 39432
rect 26283 39392 28540 39420
rect 26283 39389 26295 39392
rect 26237 39383 26295 39389
rect 28534 39380 28540 39392
rect 28592 39380 28598 39432
rect 28736 39429 28764 39460
rect 28629 39423 28687 39429
rect 28629 39389 28641 39423
rect 28675 39389 28687 39423
rect 28629 39383 28687 39389
rect 28721 39423 28779 39429
rect 28721 39389 28733 39423
rect 28767 39389 28779 39423
rect 28721 39383 28779 39389
rect 28813 39423 28871 39429
rect 28813 39389 28825 39423
rect 28859 39420 28871 39423
rect 28859 39392 28948 39420
rect 28859 39389 28871 39392
rect 28813 39383 28871 39389
rect 23750 39312 23756 39364
rect 23808 39352 23814 39364
rect 23808 39324 24532 39352
rect 23808 39312 23814 39324
rect 23014 39284 23020 39296
rect 18840 39256 23020 39284
rect 18840 39244 18846 39256
rect 23014 39244 23020 39256
rect 23072 39244 23078 39296
rect 24026 39244 24032 39296
rect 24084 39284 24090 39296
rect 24397 39287 24455 39293
rect 24397 39284 24409 39287
rect 24084 39256 24409 39284
rect 24084 39244 24090 39256
rect 24397 39253 24409 39256
rect 24443 39253 24455 39287
rect 24504 39284 24532 39324
rect 24670 39312 24676 39364
rect 24728 39352 24734 39364
rect 24857 39355 24915 39361
rect 24857 39352 24869 39355
rect 24728 39324 24869 39352
rect 24728 39312 24734 39324
rect 24857 39321 24869 39324
rect 24903 39321 24915 39355
rect 24857 39315 24915 39321
rect 25682 39312 25688 39364
rect 25740 39352 25746 39364
rect 26482 39355 26540 39361
rect 26482 39352 26494 39355
rect 25740 39324 26494 39352
rect 25740 39312 25746 39324
rect 26482 39321 26494 39324
rect 26528 39321 26540 39355
rect 26482 39315 26540 39321
rect 25130 39284 25136 39296
rect 24504 39256 25136 39284
rect 24397 39247 24455 39253
rect 25130 39244 25136 39256
rect 25188 39244 25194 39296
rect 25774 39244 25780 39296
rect 25832 39284 25838 39296
rect 27617 39287 27675 39293
rect 27617 39284 27629 39287
rect 25832 39256 27629 39284
rect 25832 39244 25838 39256
rect 27617 39253 27629 39256
rect 27663 39284 27675 39287
rect 27798 39284 27804 39296
rect 27663 39256 27804 39284
rect 27663 39253 27675 39256
rect 27617 39247 27675 39253
rect 27798 39244 27804 39256
rect 27856 39244 27862 39296
rect 28350 39284 28356 39296
rect 28311 39256 28356 39284
rect 28350 39244 28356 39256
rect 28408 39244 28414 39296
rect 28644 39284 28672 39383
rect 28920 39364 28948 39392
rect 28994 39380 29000 39432
rect 29052 39420 29058 39432
rect 29196 39420 29224 39528
rect 46290 39488 46296 39500
rect 46251 39460 46296 39488
rect 46290 39448 46296 39460
rect 46348 39448 46354 39500
rect 46477 39491 46535 39497
rect 46477 39457 46489 39491
rect 46523 39488 46535 39491
rect 47670 39488 47676 39500
rect 46523 39460 47676 39488
rect 46523 39457 46535 39460
rect 46477 39451 46535 39457
rect 47670 39448 47676 39460
rect 47728 39448 47734 39500
rect 48130 39488 48136 39500
rect 48091 39460 48136 39488
rect 48130 39448 48136 39460
rect 48188 39448 48194 39500
rect 29549 39423 29607 39429
rect 29549 39420 29561 39423
rect 29052 39392 29097 39420
rect 29196 39392 29561 39420
rect 29052 39380 29058 39392
rect 29549 39389 29561 39392
rect 29595 39389 29607 39423
rect 29549 39383 29607 39389
rect 28902 39312 28908 39364
rect 28960 39312 28966 39364
rect 28810 39284 28816 39296
rect 28644 39256 28816 39284
rect 28810 39244 28816 39256
rect 28868 39244 28874 39296
rect 29733 39287 29791 39293
rect 29733 39253 29745 39287
rect 29779 39284 29791 39287
rect 29822 39284 29828 39296
rect 29779 39256 29828 39284
rect 29779 39253 29791 39256
rect 29733 39247 29791 39253
rect 29822 39244 29828 39256
rect 29880 39244 29886 39296
rect 1104 39194 48852 39216
rect 1104 39142 19574 39194
rect 19626 39142 19638 39194
rect 19690 39142 19702 39194
rect 19754 39142 19766 39194
rect 19818 39142 19830 39194
rect 19882 39142 48852 39194
rect 1104 39120 48852 39142
rect 17402 39080 17408 39092
rect 17363 39052 17408 39080
rect 17402 39040 17408 39052
rect 17460 39040 17466 39092
rect 19797 39083 19855 39089
rect 19797 39049 19809 39083
rect 19843 39080 19855 39083
rect 20714 39080 20720 39092
rect 19843 39052 20720 39080
rect 19843 39049 19855 39052
rect 19797 39043 19855 39049
rect 20714 39040 20720 39052
rect 20772 39040 20778 39092
rect 22925 39083 22983 39089
rect 22925 39049 22937 39083
rect 22971 39080 22983 39083
rect 23842 39080 23848 39092
rect 22971 39052 23848 39080
rect 22971 39049 22983 39052
rect 22925 39043 22983 39049
rect 23842 39040 23848 39052
rect 23900 39040 23906 39092
rect 24397 39083 24455 39089
rect 24397 39049 24409 39083
rect 24443 39080 24455 39083
rect 25038 39080 25044 39092
rect 24443 39052 25044 39080
rect 24443 39049 24455 39052
rect 24397 39043 24455 39049
rect 25038 39040 25044 39052
rect 25096 39040 25102 39092
rect 25682 39080 25688 39092
rect 25643 39052 25688 39080
rect 25682 39040 25688 39052
rect 25740 39040 25746 39092
rect 27798 39080 27804 39092
rect 27759 39052 27804 39080
rect 27798 39040 27804 39052
rect 27856 39040 27862 39092
rect 29917 39083 29975 39089
rect 29917 39080 29929 39083
rect 27908 39052 29929 39080
rect 19429 39015 19487 39021
rect 19429 39012 19441 39015
rect 17880 38984 19441 39012
rect 17586 38904 17592 38956
rect 17644 38944 17650 38956
rect 17880 38953 17908 38984
rect 19429 38981 19441 38984
rect 19475 38981 19487 39015
rect 19429 38975 19487 38981
rect 19702 38972 19708 39024
rect 19760 39012 19766 39024
rect 22833 39015 22891 39021
rect 22833 39012 22845 39015
rect 19760 38984 22845 39012
rect 19760 38972 19766 38984
rect 22833 38981 22845 38984
rect 22879 38981 22891 39015
rect 24026 39012 24032 39024
rect 23987 38984 24032 39012
rect 22833 38975 22891 38981
rect 24026 38972 24032 38984
rect 24084 38972 24090 39024
rect 24946 39012 24952 39024
rect 24136 38984 24952 39012
rect 17681 38947 17739 38953
rect 17681 38944 17693 38947
rect 17644 38916 17693 38944
rect 17644 38904 17650 38916
rect 17681 38913 17693 38916
rect 17727 38913 17739 38947
rect 17681 38907 17739 38913
rect 17773 38947 17831 38953
rect 17773 38913 17785 38947
rect 17819 38913 17831 38947
rect 17773 38907 17831 38913
rect 17865 38947 17923 38953
rect 17865 38913 17877 38947
rect 17911 38913 17923 38947
rect 17865 38907 17923 38913
rect 18049 38947 18107 38953
rect 18049 38913 18061 38947
rect 18095 38913 18107 38947
rect 18506 38944 18512 38956
rect 18467 38916 18512 38944
rect 18049 38907 18107 38913
rect 2038 38876 2044 38888
rect 1999 38848 2044 38876
rect 2038 38836 2044 38848
rect 2096 38836 2102 38888
rect 2225 38879 2283 38885
rect 2225 38845 2237 38879
rect 2271 38876 2283 38879
rect 2774 38876 2780 38888
rect 2271 38848 2780 38876
rect 2271 38845 2283 38848
rect 2225 38839 2283 38845
rect 2774 38836 2780 38848
rect 2832 38836 2838 38888
rect 2866 38836 2872 38888
rect 2924 38876 2930 38888
rect 2924 38848 2969 38876
rect 2924 38836 2930 38848
rect 17788 38740 17816 38907
rect 17862 38768 17868 38820
rect 17920 38808 17926 38820
rect 18064 38808 18092 38907
rect 18506 38904 18512 38916
rect 18564 38904 18570 38956
rect 19613 38947 19671 38953
rect 19613 38913 19625 38947
rect 19659 38944 19671 38947
rect 19794 38944 19800 38956
rect 19659 38916 19800 38944
rect 19659 38913 19671 38916
rect 19613 38907 19671 38913
rect 19794 38904 19800 38916
rect 19852 38904 19858 38956
rect 19889 38947 19947 38953
rect 19889 38913 19901 38947
rect 19935 38944 19947 38947
rect 24136 38944 24164 38984
rect 24946 38972 24952 38984
rect 25004 38972 25010 39024
rect 25130 38972 25136 39024
rect 25188 39012 25194 39024
rect 25188 38984 26372 39012
rect 25188 38972 25194 38984
rect 19935 38916 24164 38944
rect 19935 38913 19947 38916
rect 19889 38907 19947 38913
rect 18690 38836 18696 38888
rect 18748 38876 18754 38888
rect 19904 38876 19932 38907
rect 24210 38904 24216 38956
rect 24268 38944 24274 38956
rect 24857 38947 24915 38953
rect 24268 38916 24313 38944
rect 24268 38904 24274 38916
rect 24857 38913 24869 38947
rect 24903 38944 24915 38947
rect 25774 38944 25780 38956
rect 24903 38916 25780 38944
rect 24903 38913 24915 38916
rect 24857 38907 24915 38913
rect 25774 38904 25780 38916
rect 25832 38904 25838 38956
rect 25961 38947 26019 38953
rect 25961 38913 25973 38947
rect 26007 38913 26019 38947
rect 25961 38907 26019 38913
rect 26053 38947 26111 38953
rect 26053 38913 26065 38947
rect 26099 38913 26111 38947
rect 26053 38907 26111 38913
rect 18748 38848 19932 38876
rect 18748 38836 18754 38848
rect 22278 38836 22284 38888
rect 22336 38876 22342 38888
rect 24949 38879 25007 38885
rect 24949 38876 24961 38879
rect 22336 38848 24961 38876
rect 22336 38836 22342 38848
rect 24949 38845 24961 38848
rect 24995 38845 25007 38879
rect 24949 38839 25007 38845
rect 25222 38836 25228 38888
rect 25280 38876 25286 38888
rect 25976 38876 26004 38907
rect 25280 38848 26004 38876
rect 25280 38836 25286 38848
rect 26068 38808 26096 38907
rect 26142 38904 26148 38956
rect 26200 38944 26206 38956
rect 26344 38953 26372 38984
rect 27338 38972 27344 39024
rect 27396 39012 27402 39024
rect 27908 39012 27936 39052
rect 29917 39049 29929 39052
rect 29963 39049 29975 39083
rect 48038 39080 48044 39092
rect 47999 39052 48044 39080
rect 29917 39043 29975 39049
rect 48038 39040 48044 39052
rect 48096 39040 48102 39092
rect 27396 38984 27936 39012
rect 27396 38972 27402 38984
rect 28350 38972 28356 39024
rect 28408 39012 28414 39024
rect 28782 39015 28840 39021
rect 28782 39012 28794 39015
rect 28408 38984 28794 39012
rect 28408 38972 28414 38984
rect 28782 38981 28794 38984
rect 28828 38981 28840 39015
rect 28782 38975 28840 38981
rect 26329 38947 26387 38953
rect 26200 38916 26245 38944
rect 26200 38904 26206 38916
rect 26329 38913 26341 38947
rect 26375 38913 26387 38947
rect 26329 38907 26387 38913
rect 27709 38947 27767 38953
rect 27709 38913 27721 38947
rect 27755 38944 27767 38947
rect 27798 38944 27804 38956
rect 27755 38916 27804 38944
rect 27755 38913 27767 38916
rect 27709 38907 27767 38913
rect 27798 38904 27804 38916
rect 27856 38904 27862 38956
rect 28534 38944 28540 38956
rect 28495 38916 28540 38944
rect 28534 38904 28540 38916
rect 28592 38904 28598 38956
rect 47946 38944 47952 38956
rect 47907 38916 47952 38944
rect 47946 38904 47952 38916
rect 48004 38904 48010 38956
rect 27522 38876 27528 38888
rect 17920 38780 18092 38808
rect 24044 38780 26096 38808
rect 26712 38848 27528 38876
rect 17920 38768 17926 38780
rect 18693 38743 18751 38749
rect 18693 38740 18705 38743
rect 17788 38712 18705 38740
rect 18693 38709 18705 38712
rect 18739 38740 18751 38743
rect 18782 38740 18788 38752
rect 18739 38712 18788 38740
rect 18739 38709 18751 38712
rect 18693 38703 18751 38709
rect 18782 38700 18788 38712
rect 18840 38740 18846 38752
rect 24044 38740 24072 38780
rect 24946 38740 24952 38752
rect 18840 38712 24072 38740
rect 24907 38712 24952 38740
rect 18840 38700 18846 38712
rect 24946 38700 24952 38712
rect 25004 38700 25010 38752
rect 25130 38700 25136 38752
rect 25188 38740 25194 38752
rect 25225 38743 25283 38749
rect 25225 38740 25237 38743
rect 25188 38712 25237 38740
rect 25188 38700 25194 38712
rect 25225 38709 25237 38712
rect 25271 38709 25283 38743
rect 25225 38703 25283 38709
rect 26050 38700 26056 38752
rect 26108 38740 26114 38752
rect 26712 38740 26740 38848
rect 27522 38836 27528 38848
rect 27580 38876 27586 38888
rect 27893 38879 27951 38885
rect 27893 38876 27905 38879
rect 27580 38848 27905 38876
rect 27580 38836 27586 38848
rect 27893 38845 27905 38848
rect 27939 38845 27951 38879
rect 27893 38839 27951 38845
rect 27338 38740 27344 38752
rect 26108 38712 26740 38740
rect 27299 38712 27344 38740
rect 26108 38700 26114 38712
rect 27338 38700 27344 38712
rect 27396 38700 27402 38752
rect 47026 38740 47032 38752
rect 46987 38712 47032 38740
rect 47026 38700 47032 38712
rect 47084 38700 47090 38752
rect 1104 38650 48852 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 48852 38650
rect 1104 38576 48852 38598
rect 2038 38496 2044 38548
rect 2096 38536 2102 38548
rect 2317 38539 2375 38545
rect 2317 38536 2329 38539
rect 2096 38508 2329 38536
rect 2096 38496 2102 38508
rect 2317 38505 2329 38508
rect 2363 38505 2375 38539
rect 2317 38499 2375 38505
rect 21266 38496 21272 38548
rect 21324 38536 21330 38548
rect 22922 38536 22928 38548
rect 21324 38508 22928 38536
rect 21324 38496 21330 38508
rect 22922 38496 22928 38508
rect 22980 38536 22986 38548
rect 23109 38539 23167 38545
rect 23109 38536 23121 38539
rect 22980 38508 23121 38536
rect 22980 38496 22986 38508
rect 23109 38505 23121 38508
rect 23155 38505 23167 38539
rect 23109 38499 23167 38505
rect 23569 38539 23627 38545
rect 23569 38505 23581 38539
rect 23615 38536 23627 38539
rect 24949 38539 25007 38545
rect 24949 38536 24961 38539
rect 23615 38508 24961 38536
rect 23615 38505 23627 38508
rect 23569 38499 23627 38505
rect 24949 38505 24961 38508
rect 24995 38505 25007 38539
rect 24949 38499 25007 38505
rect 27798 38496 27804 38548
rect 27856 38536 27862 38548
rect 30929 38539 30987 38545
rect 30929 38536 30941 38539
rect 27856 38508 30941 38536
rect 27856 38496 27862 38508
rect 30929 38505 30941 38508
rect 30975 38505 30987 38539
rect 30929 38499 30987 38505
rect 17773 38471 17831 38477
rect 17773 38437 17785 38471
rect 17819 38468 17831 38471
rect 17862 38468 17868 38480
rect 17819 38440 17868 38468
rect 17819 38437 17831 38440
rect 17773 38431 17831 38437
rect 17862 38428 17868 38440
rect 17920 38428 17926 38480
rect 19889 38471 19947 38477
rect 19889 38437 19901 38471
rect 19935 38468 19947 38471
rect 20070 38468 20076 38480
rect 19935 38440 20076 38468
rect 19935 38437 19947 38440
rect 19889 38431 19947 38437
rect 20070 38428 20076 38440
rect 20128 38428 20134 38480
rect 25314 38468 25320 38480
rect 20180 38440 25320 38468
rect 18414 38360 18420 38412
rect 18472 38400 18478 38412
rect 20180 38400 20208 38440
rect 25314 38428 25320 38440
rect 25372 38428 25378 38480
rect 28534 38428 28540 38480
rect 28592 38468 28598 38480
rect 28592 38440 29592 38468
rect 28592 38428 28598 38440
rect 18472 38372 20208 38400
rect 18472 38360 18478 38372
rect 22094 38360 22100 38412
rect 22152 38400 22158 38412
rect 23106 38400 23112 38412
rect 22152 38372 23112 38400
rect 22152 38360 22158 38372
rect 23106 38360 23112 38372
rect 23164 38400 23170 38412
rect 23201 38403 23259 38409
rect 23201 38400 23213 38403
rect 23164 38372 23213 38400
rect 23164 38360 23170 38372
rect 23201 38369 23213 38372
rect 23247 38369 23259 38403
rect 23201 38363 23259 38369
rect 24210 38360 24216 38412
rect 24268 38400 24274 38412
rect 28074 38400 28080 38412
rect 24268 38372 28080 38400
rect 24268 38360 24274 38372
rect 17589 38335 17647 38341
rect 17589 38301 17601 38335
rect 17635 38332 17647 38335
rect 17635 38304 19380 38332
rect 17635 38301 17647 38304
rect 17589 38295 17647 38301
rect 19352 38276 19380 38304
rect 21082 38292 21088 38344
rect 21140 38332 21146 38344
rect 22235 38335 22293 38341
rect 22235 38332 22247 38335
rect 21140 38304 22247 38332
rect 21140 38292 21146 38304
rect 22235 38301 22247 38304
rect 22281 38301 22293 38335
rect 22370 38332 22376 38344
rect 22331 38304 22376 38332
rect 22235 38295 22293 38301
rect 22370 38292 22376 38304
rect 22428 38292 22434 38344
rect 22480 38341 22600 38342
rect 22465 38335 22600 38341
rect 22465 38301 22477 38335
rect 22511 38314 22600 38335
rect 22511 38301 22523 38314
rect 22465 38295 22523 38301
rect 17034 38224 17040 38276
rect 17092 38264 17098 38276
rect 18325 38267 18383 38273
rect 18325 38264 18337 38267
rect 17092 38236 18337 38264
rect 17092 38224 17098 38236
rect 18325 38233 18337 38236
rect 18371 38264 18383 38267
rect 18506 38264 18512 38276
rect 18371 38236 18512 38264
rect 18371 38233 18383 38236
rect 18325 38227 18383 38233
rect 18506 38224 18512 38236
rect 18564 38224 18570 38276
rect 19334 38224 19340 38276
rect 19392 38264 19398 38276
rect 19702 38264 19708 38276
rect 19392 38236 19708 38264
rect 19392 38224 19398 38236
rect 19702 38224 19708 38236
rect 19760 38224 19766 38276
rect 22572 38264 22600 38314
rect 22649 38335 22707 38341
rect 22649 38301 22661 38335
rect 22695 38332 22707 38335
rect 22830 38332 22836 38344
rect 22695 38304 22836 38332
rect 22695 38301 22707 38304
rect 22649 38295 22707 38301
rect 22830 38292 22836 38304
rect 22888 38292 22894 38344
rect 23385 38335 23443 38341
rect 23385 38301 23397 38335
rect 23431 38332 23443 38335
rect 23566 38332 23572 38344
rect 23431 38304 23572 38332
rect 23431 38301 23443 38304
rect 23385 38295 23443 38301
rect 23566 38292 23572 38304
rect 23624 38292 23630 38344
rect 24946 38332 24952 38344
rect 24907 38304 24952 38332
rect 24946 38292 24952 38304
rect 25004 38292 25010 38344
rect 25130 38332 25136 38344
rect 25091 38304 25136 38332
rect 25130 38292 25136 38304
rect 25188 38292 25194 38344
rect 27338 38292 27344 38344
rect 27396 38332 27402 38344
rect 27724 38341 27752 38372
rect 28074 38360 28080 38372
rect 28132 38360 28138 38412
rect 28442 38360 28448 38412
rect 28500 38400 28506 38412
rect 29564 38409 29592 38440
rect 29549 38403 29607 38409
rect 28500 38372 28764 38400
rect 28500 38360 28506 38372
rect 27525 38335 27583 38341
rect 27525 38332 27537 38335
rect 27396 38304 27537 38332
rect 27396 38292 27402 38304
rect 27525 38301 27537 38304
rect 27571 38301 27583 38335
rect 27525 38295 27583 38301
rect 27709 38335 27767 38341
rect 27709 38301 27721 38335
rect 27755 38301 27767 38335
rect 28626 38332 28632 38344
rect 28587 38304 28632 38332
rect 27709 38295 27767 38301
rect 28626 38292 28632 38304
rect 28684 38292 28690 38344
rect 28736 38341 28764 38372
rect 29549 38369 29561 38403
rect 29595 38369 29607 38403
rect 29549 38363 29607 38369
rect 46293 38403 46351 38409
rect 46293 38369 46305 38403
rect 46339 38400 46351 38403
rect 47026 38400 47032 38412
rect 46339 38372 47032 38400
rect 46339 38369 46351 38372
rect 46293 38363 46351 38369
rect 47026 38360 47032 38372
rect 47084 38360 47090 38412
rect 48133 38403 48191 38409
rect 48133 38369 48145 38403
rect 48179 38400 48191 38403
rect 48222 38400 48228 38412
rect 48179 38372 48228 38400
rect 48179 38369 48191 38372
rect 48133 38363 48191 38369
rect 48222 38360 48228 38372
rect 48280 38360 48286 38412
rect 28721 38335 28779 38341
rect 28721 38301 28733 38335
rect 28767 38301 28779 38335
rect 28721 38295 28779 38301
rect 28813 38335 28871 38341
rect 28813 38301 28825 38335
rect 28859 38332 28871 38335
rect 28902 38332 28908 38344
rect 28859 38304 28908 38332
rect 28859 38301 28871 38304
rect 28813 38295 28871 38301
rect 28902 38292 28908 38304
rect 28960 38292 28966 38344
rect 28997 38335 29055 38341
rect 28997 38301 29009 38335
rect 29043 38332 29055 38335
rect 29086 38332 29092 38344
rect 29043 38304 29092 38332
rect 29043 38301 29055 38304
rect 28997 38295 29055 38301
rect 29086 38292 29092 38304
rect 29144 38292 29150 38344
rect 23014 38264 23020 38276
rect 22572 38236 23020 38264
rect 23014 38224 23020 38236
rect 23072 38224 23078 38276
rect 23109 38267 23167 38273
rect 23109 38233 23121 38267
rect 23155 38264 23167 38267
rect 24670 38264 24676 38276
rect 23155 38236 24676 38264
rect 23155 38233 23167 38236
rect 23109 38227 23167 38233
rect 24670 38224 24676 38236
rect 24728 38224 24734 38276
rect 28353 38267 28411 38273
rect 28353 38233 28365 38267
rect 28399 38264 28411 38267
rect 29794 38267 29852 38273
rect 29794 38264 29806 38267
rect 28399 38236 29806 38264
rect 28399 38233 28411 38236
rect 28353 38227 28411 38233
rect 29794 38233 29806 38236
rect 29840 38233 29852 38267
rect 29794 38227 29852 38233
rect 46477 38267 46535 38273
rect 46477 38233 46489 38267
rect 46523 38264 46535 38267
rect 46934 38264 46940 38276
rect 46523 38236 46940 38264
rect 46523 38233 46535 38236
rect 46477 38227 46535 38233
rect 46934 38224 46940 38236
rect 46992 38224 46998 38276
rect 18414 38196 18420 38208
rect 18375 38168 18420 38196
rect 18414 38156 18420 38168
rect 18472 38156 18478 38208
rect 22002 38196 22008 38208
rect 21963 38168 22008 38196
rect 22002 38156 22008 38168
rect 22060 38156 22066 38208
rect 25317 38199 25375 38205
rect 25317 38165 25329 38199
rect 25363 38196 25375 38199
rect 25682 38196 25688 38208
rect 25363 38168 25688 38196
rect 25363 38165 25375 38168
rect 25317 38159 25375 38165
rect 25682 38156 25688 38168
rect 25740 38156 25746 38208
rect 27893 38199 27951 38205
rect 27893 38165 27905 38199
rect 27939 38196 27951 38199
rect 28902 38196 28908 38208
rect 27939 38168 28908 38196
rect 27939 38165 27951 38168
rect 27893 38159 27951 38165
rect 28902 38156 28908 38168
rect 28960 38156 28966 38208
rect 1104 38106 48852 38128
rect 1104 38054 19574 38106
rect 19626 38054 19638 38106
rect 19690 38054 19702 38106
rect 19754 38054 19766 38106
rect 19818 38054 19830 38106
rect 19882 38054 48852 38106
rect 1104 38032 48852 38054
rect 2774 37952 2780 38004
rect 2832 37992 2838 38004
rect 3053 37995 3111 38001
rect 3053 37992 3065 37995
rect 2832 37964 3065 37992
rect 2832 37952 2838 37964
rect 3053 37961 3065 37964
rect 3099 37961 3111 37995
rect 3053 37955 3111 37961
rect 23845 37995 23903 38001
rect 23845 37961 23857 37995
rect 23891 37992 23903 37995
rect 24673 37995 24731 38001
rect 24673 37992 24685 37995
rect 23891 37964 24685 37992
rect 23891 37961 23903 37964
rect 23845 37955 23903 37961
rect 24673 37961 24685 37964
rect 24719 37992 24731 37995
rect 24854 37992 24860 38004
rect 24719 37964 24860 37992
rect 24719 37961 24731 37964
rect 24673 37955 24731 37961
rect 24854 37952 24860 37964
rect 24912 37952 24918 38004
rect 24946 37952 24952 38004
rect 25004 37992 25010 38004
rect 25961 37995 26019 38001
rect 25961 37992 25973 37995
rect 25004 37964 25973 37992
rect 25004 37952 25010 37964
rect 25961 37961 25973 37964
rect 26007 37961 26019 37995
rect 46934 37992 46940 38004
rect 46895 37964 46940 37992
rect 25961 37955 26019 37961
rect 46934 37952 46940 37964
rect 46992 37952 46998 38004
rect 17126 37884 17132 37936
rect 17184 37924 17190 37936
rect 17184 37896 20116 37924
rect 17184 37884 17190 37896
rect 1854 37856 1860 37868
rect 1815 37828 1860 37856
rect 1854 37816 1860 37828
rect 1912 37816 1918 37868
rect 2961 37859 3019 37865
rect 2961 37825 2973 37859
rect 3007 37856 3019 37859
rect 7282 37856 7288 37868
rect 3007 37828 7288 37856
rect 3007 37825 3019 37828
rect 2961 37819 3019 37825
rect 7282 37816 7288 37828
rect 7340 37816 7346 37868
rect 18233 37859 18291 37865
rect 18233 37825 18245 37859
rect 18279 37856 18291 37859
rect 18322 37856 18328 37868
rect 18279 37828 18328 37856
rect 18279 37825 18291 37828
rect 18233 37819 18291 37825
rect 18322 37816 18328 37828
rect 18380 37816 18386 37868
rect 18417 37859 18475 37865
rect 18417 37825 18429 37859
rect 18463 37856 18475 37859
rect 19426 37856 19432 37868
rect 18463 37828 19432 37856
rect 18463 37825 18475 37828
rect 18417 37819 18475 37825
rect 19426 37816 19432 37828
rect 19484 37816 19490 37868
rect 20088 37856 20116 37896
rect 22002 37884 22008 37936
rect 22060 37924 22066 37936
rect 22710 37927 22768 37933
rect 22710 37924 22722 37927
rect 22060 37896 22722 37924
rect 22060 37884 22066 37896
rect 22710 37893 22722 37896
rect 22756 37893 22768 37927
rect 22710 37887 22768 37893
rect 22830 37884 22836 37936
rect 22888 37884 22894 37936
rect 24765 37927 24823 37933
rect 24765 37893 24777 37927
rect 24811 37924 24823 37927
rect 24811 37896 25636 37924
rect 24811 37893 24823 37896
rect 24765 37887 24823 37893
rect 20855 37859 20913 37865
rect 20855 37856 20867 37859
rect 20088 37828 20867 37856
rect 20855 37825 20867 37828
rect 20901 37825 20913 37859
rect 20855 37819 20913 37825
rect 20974 37862 21032 37868
rect 20974 37828 20986 37862
rect 21020 37828 21032 37862
rect 20974 37822 21032 37828
rect 21090 37859 21148 37865
rect 21090 37825 21102 37859
rect 21136 37825 21148 37859
rect 20989 37732 21017 37822
rect 21090 37819 21148 37825
rect 21269 37859 21327 37865
rect 21269 37825 21281 37859
rect 21315 37856 21327 37859
rect 22370 37856 22376 37868
rect 21315 37828 22376 37856
rect 21315 37825 21327 37828
rect 21269 37819 21327 37825
rect 21100 37788 21128 37819
rect 22370 37816 22376 37828
rect 22428 37856 22434 37868
rect 22848 37856 22876 37884
rect 22428 37828 22876 37856
rect 22428 37816 22434 37828
rect 25130 37816 25136 37868
rect 25188 37856 25194 37868
rect 25501 37859 25559 37865
rect 25501 37856 25513 37859
rect 25188 37828 25513 37856
rect 25188 37816 25194 37828
rect 25501 37825 25513 37828
rect 25547 37825 25559 37859
rect 25501 37819 25559 37825
rect 21174 37788 21180 37800
rect 21100 37760 21180 37788
rect 21174 37748 21180 37760
rect 21232 37748 21238 37800
rect 22186 37748 22192 37800
rect 22244 37788 22250 37800
rect 22465 37791 22523 37797
rect 22465 37788 22477 37791
rect 22244 37760 22477 37788
rect 22244 37748 22250 37760
rect 22465 37757 22477 37760
rect 22511 37757 22523 37791
rect 24946 37788 24952 37800
rect 24907 37760 24952 37788
rect 22465 37751 22523 37757
rect 24946 37748 24952 37760
rect 25004 37748 25010 37800
rect 25608 37788 25636 37896
rect 28994 37884 29000 37936
rect 29052 37924 29058 37936
rect 29052 37896 29592 37924
rect 29052 37884 29058 37896
rect 25774 37856 25780 37868
rect 25735 37828 25780 37856
rect 25774 37816 25780 37828
rect 25832 37816 25838 37868
rect 29178 37856 29184 37868
rect 29139 37828 29184 37856
rect 29178 37816 29184 37828
rect 29236 37816 29242 37868
rect 29273 37859 29331 37865
rect 29273 37825 29285 37859
rect 29319 37825 29331 37859
rect 29273 37819 29331 37825
rect 25685 37791 25743 37797
rect 25685 37788 25697 37791
rect 25608 37760 25697 37788
rect 25685 37757 25697 37760
rect 25731 37788 25743 37791
rect 27798 37788 27804 37800
rect 25731 37760 27804 37788
rect 25731 37757 25743 37760
rect 25685 37751 25743 37757
rect 27798 37748 27804 37760
rect 27856 37748 27862 37800
rect 20989 37692 20996 37732
rect 20990 37680 20996 37692
rect 21048 37680 21054 37732
rect 25314 37680 25320 37732
rect 25372 37720 25378 37732
rect 28442 37720 28448 37732
rect 25372 37692 28448 37720
rect 25372 37680 25378 37692
rect 28442 37680 28448 37692
rect 28500 37720 28506 37732
rect 29288 37720 29316 37819
rect 29362 37816 29368 37868
rect 29420 37856 29426 37868
rect 29564 37865 29592 37896
rect 29549 37859 29607 37865
rect 29420 37828 29465 37856
rect 29420 37816 29426 37828
rect 29549 37825 29561 37859
rect 29595 37825 29607 37859
rect 29549 37819 29607 37825
rect 46845 37859 46903 37865
rect 46845 37825 46857 37859
rect 46891 37856 46903 37859
rect 47302 37856 47308 37868
rect 46891 37828 47308 37856
rect 46891 37825 46903 37828
rect 46845 37819 46903 37825
rect 47302 37816 47308 37828
rect 47360 37816 47366 37868
rect 47854 37856 47860 37868
rect 47815 37828 47860 37856
rect 47854 37816 47860 37828
rect 47912 37816 47918 37868
rect 28500 37692 29316 37720
rect 28500 37680 28506 37692
rect 1946 37652 1952 37664
rect 1907 37624 1952 37652
rect 1946 37612 1952 37624
rect 2004 37612 2010 37664
rect 18598 37652 18604 37664
rect 18559 37624 18604 37652
rect 18598 37612 18604 37624
rect 18656 37612 18662 37664
rect 20625 37655 20683 37661
rect 20625 37621 20637 37655
rect 20671 37652 20683 37655
rect 21082 37652 21088 37664
rect 20671 37624 21088 37652
rect 20671 37621 20683 37624
rect 20625 37615 20683 37621
rect 21082 37612 21088 37624
rect 21140 37612 21146 37664
rect 24302 37652 24308 37664
rect 24263 37624 24308 37652
rect 24302 37612 24308 37624
rect 24360 37612 24366 37664
rect 25777 37655 25835 37661
rect 25777 37621 25789 37655
rect 25823 37652 25835 37655
rect 26234 37652 26240 37664
rect 25823 37624 26240 37652
rect 25823 37621 25835 37624
rect 25777 37615 25835 37621
rect 26234 37612 26240 37624
rect 26292 37652 26298 37664
rect 27246 37652 27252 37664
rect 26292 37624 27252 37652
rect 26292 37612 26298 37624
rect 27246 37612 27252 37624
rect 27304 37612 27310 37664
rect 28905 37655 28963 37661
rect 28905 37621 28917 37655
rect 28951 37652 28963 37655
rect 29638 37652 29644 37664
rect 28951 37624 29644 37652
rect 28951 37621 28963 37624
rect 28905 37615 28963 37621
rect 29638 37612 29644 37624
rect 29696 37612 29702 37664
rect 48038 37652 48044 37664
rect 47999 37624 48044 37652
rect 48038 37612 48044 37624
rect 48096 37612 48102 37664
rect 1104 37562 48852 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 48852 37562
rect 1104 37488 48852 37510
rect 1946 37408 1952 37460
rect 2004 37448 2010 37460
rect 2004 37420 18276 37448
rect 2004 37408 2010 37420
rect 18248 37380 18276 37420
rect 18322 37408 18328 37460
rect 18380 37448 18386 37460
rect 19245 37451 19303 37457
rect 19245 37448 19257 37451
rect 18380 37420 19257 37448
rect 18380 37408 18386 37420
rect 19245 37417 19257 37420
rect 19291 37417 19303 37451
rect 19245 37411 19303 37417
rect 23014 37408 23020 37460
rect 23072 37448 23078 37460
rect 23845 37451 23903 37457
rect 23845 37448 23857 37451
rect 23072 37420 23857 37448
rect 23072 37408 23078 37420
rect 23845 37417 23857 37420
rect 23891 37417 23903 37451
rect 23845 37411 23903 37417
rect 19150 37380 19156 37392
rect 18248 37352 19156 37380
rect 19150 37340 19156 37352
rect 19208 37340 19214 37392
rect 26234 37380 26240 37392
rect 24872 37352 26240 37380
rect 1394 37312 1400 37324
rect 1355 37284 1400 37312
rect 1394 37272 1400 37284
rect 1452 37272 1458 37324
rect 4062 37272 4068 37324
rect 4120 37312 4126 37324
rect 8294 37312 8300 37324
rect 4120 37284 8300 37312
rect 4120 37272 4126 37284
rect 8294 37272 8300 37284
rect 8352 37272 8358 37324
rect 19058 37272 19064 37324
rect 19116 37312 19122 37324
rect 19334 37312 19340 37324
rect 19116 37284 19340 37312
rect 19116 37272 19122 37284
rect 19334 37272 19340 37284
rect 19392 37272 19398 37324
rect 19889 37315 19947 37321
rect 19889 37281 19901 37315
rect 19935 37312 19947 37315
rect 19978 37312 19984 37324
rect 19935 37284 19984 37312
rect 19935 37281 19947 37284
rect 19889 37275 19947 37281
rect 19978 37272 19984 37284
rect 20036 37272 20042 37324
rect 22738 37272 22744 37324
rect 22796 37312 22802 37324
rect 24872 37321 24900 37352
rect 26234 37340 26240 37352
rect 26292 37340 26298 37392
rect 27798 37340 27804 37392
rect 27856 37380 27862 37392
rect 27893 37383 27951 37389
rect 27893 37380 27905 37383
rect 27856 37352 27905 37380
rect 27856 37340 27862 37352
rect 27893 37349 27905 37352
rect 27939 37380 27951 37383
rect 28534 37380 28540 37392
rect 27939 37352 28540 37380
rect 27939 37349 27951 37352
rect 27893 37343 27951 37349
rect 28534 37340 28540 37352
rect 28592 37380 28598 37392
rect 28592 37352 29592 37380
rect 28592 37340 28598 37352
rect 24857 37315 24915 37321
rect 22796 37284 24808 37312
rect 22796 37272 22802 37284
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37244 1731 37247
rect 7282 37244 7288 37256
rect 1719 37216 2774 37244
rect 7243 37216 7288 37244
rect 1719 37213 1731 37216
rect 1673 37207 1731 37213
rect 2130 37136 2136 37188
rect 2188 37176 2194 37188
rect 2314 37176 2320 37188
rect 2188 37148 2320 37176
rect 2188 37136 2194 37148
rect 2314 37136 2320 37148
rect 2372 37136 2378 37188
rect 2746 37176 2774 37216
rect 7282 37204 7288 37216
rect 7340 37204 7346 37256
rect 16482 37204 16488 37256
rect 16540 37244 16546 37256
rect 17313 37247 17371 37253
rect 17313 37244 17325 37247
rect 16540 37216 17325 37244
rect 16540 37204 16546 37216
rect 17313 37213 17325 37216
rect 17359 37213 17371 37247
rect 17313 37207 17371 37213
rect 19705 37247 19763 37253
rect 19705 37213 19717 37247
rect 19751 37244 19763 37247
rect 20438 37244 20444 37256
rect 19751 37216 20444 37244
rect 19751 37213 19763 37216
rect 19705 37207 19763 37213
rect 20438 37204 20444 37216
rect 20496 37204 20502 37256
rect 20622 37204 20628 37256
rect 20680 37244 20686 37256
rect 20993 37247 21051 37253
rect 20993 37244 21005 37247
rect 20680 37216 21005 37244
rect 20680 37204 20686 37216
rect 20993 37213 21005 37216
rect 21039 37213 21051 37247
rect 20993 37207 21051 37213
rect 21082 37204 21088 37256
rect 21140 37244 21146 37256
rect 21249 37247 21307 37253
rect 21249 37244 21261 37247
rect 21140 37216 21261 37244
rect 21140 37204 21146 37216
rect 21249 37213 21261 37216
rect 21295 37213 21307 37247
rect 21249 37207 21307 37213
rect 23477 37247 23535 37253
rect 23477 37213 23489 37247
rect 23523 37244 23535 37247
rect 24302 37244 24308 37256
rect 23523 37216 24308 37244
rect 23523 37213 23535 37216
rect 23477 37207 23535 37213
rect 24302 37204 24308 37216
rect 24360 37204 24366 37256
rect 24780 37253 24808 37284
rect 24857 37281 24869 37315
rect 24903 37281 24915 37315
rect 24857 37275 24915 37281
rect 24946 37272 24952 37324
rect 25004 37312 25010 37324
rect 25041 37315 25099 37321
rect 25041 37312 25053 37315
rect 25004 37284 25053 37312
rect 25004 37272 25010 37284
rect 25041 37281 25053 37284
rect 25087 37312 25099 37315
rect 26142 37312 26148 37324
rect 25087 37284 26148 37312
rect 25087 37281 25099 37284
rect 25041 37275 25099 37281
rect 26142 37272 26148 37284
rect 26200 37272 26206 37324
rect 29564 37321 29592 37352
rect 29549 37315 29607 37321
rect 29549 37281 29561 37315
rect 29595 37281 29607 37315
rect 29549 37275 29607 37281
rect 33042 37272 33048 37324
rect 33100 37312 33106 37324
rect 46842 37312 46848 37324
rect 33100 37284 46848 37312
rect 33100 37272 33106 37284
rect 46842 37272 46848 37284
rect 46900 37272 46906 37324
rect 24765 37247 24823 37253
rect 24765 37213 24777 37247
rect 24811 37213 24823 37247
rect 24765 37207 24823 37213
rect 29638 37204 29644 37256
rect 29696 37244 29702 37256
rect 29805 37247 29863 37253
rect 29805 37244 29817 37247
rect 29696 37216 29817 37244
rect 29696 37204 29702 37216
rect 29805 37213 29817 37216
rect 29851 37213 29863 37247
rect 46290 37244 46296 37256
rect 46251 37216 46296 37244
rect 29805 37207 29863 37213
rect 46290 37204 46296 37216
rect 46348 37204 46354 37256
rect 17218 37176 17224 37188
rect 2746 37148 17224 37176
rect 17218 37136 17224 37148
rect 17276 37136 17282 37188
rect 17580 37179 17638 37185
rect 17580 37145 17592 37179
rect 17626 37176 17638 37179
rect 17678 37176 17684 37188
rect 17626 37148 17684 37176
rect 17626 37145 17638 37148
rect 17580 37139 17638 37145
rect 17678 37136 17684 37148
rect 17736 37136 17742 37188
rect 19613 37179 19671 37185
rect 19613 37176 19625 37179
rect 18708 37148 19625 37176
rect 7374 37108 7380 37120
rect 7335 37080 7380 37108
rect 7374 37068 7380 37080
rect 7432 37068 7438 37120
rect 18708 37117 18736 37148
rect 19613 37145 19625 37148
rect 19659 37176 19671 37179
rect 23661 37179 23719 37185
rect 19659 37148 23612 37176
rect 19659 37145 19671 37148
rect 19613 37139 19671 37145
rect 18693 37111 18751 37117
rect 18693 37077 18705 37111
rect 18739 37077 18751 37111
rect 18693 37071 18751 37077
rect 22373 37111 22431 37117
rect 22373 37077 22385 37111
rect 22419 37108 22431 37111
rect 22738 37108 22744 37120
rect 22419 37080 22744 37108
rect 22419 37077 22431 37080
rect 22373 37071 22431 37077
rect 22738 37068 22744 37080
rect 22796 37068 22802 37120
rect 23584 37108 23612 37148
rect 23661 37145 23673 37179
rect 23707 37176 23719 37179
rect 23750 37176 23756 37188
rect 23707 37148 23756 37176
rect 23707 37145 23719 37148
rect 23661 37139 23719 37145
rect 23750 37136 23756 37148
rect 23808 37136 23814 37188
rect 25774 37176 25780 37188
rect 24228 37148 25780 37176
rect 24228 37108 24256 37148
rect 25774 37136 25780 37148
rect 25832 37136 25838 37188
rect 27062 37136 27068 37188
rect 27120 37176 27126 37188
rect 27709 37179 27767 37185
rect 27709 37176 27721 37179
rect 27120 37148 27721 37176
rect 27120 37136 27126 37148
rect 27709 37145 27721 37148
rect 27755 37145 27767 37179
rect 27709 37139 27767 37145
rect 46477 37179 46535 37185
rect 46477 37145 46489 37179
rect 46523 37176 46535 37179
rect 47670 37176 47676 37188
rect 46523 37148 47676 37176
rect 46523 37145 46535 37148
rect 46477 37139 46535 37145
rect 47670 37136 47676 37148
rect 47728 37136 47734 37188
rect 48130 37176 48136 37188
rect 48091 37148 48136 37176
rect 48130 37136 48136 37148
rect 48188 37136 48194 37188
rect 24394 37108 24400 37120
rect 23584 37080 24256 37108
rect 24355 37080 24400 37108
rect 24394 37068 24400 37080
rect 24452 37068 24458 37120
rect 25866 37068 25872 37120
rect 25924 37108 25930 37120
rect 29638 37108 29644 37120
rect 25924 37080 29644 37108
rect 25924 37068 25930 37080
rect 29638 37068 29644 37080
rect 29696 37068 29702 37120
rect 30926 37108 30932 37120
rect 30887 37080 30932 37108
rect 30926 37068 30932 37080
rect 30984 37068 30990 37120
rect 1104 37018 48852 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 48852 37018
rect 1104 36944 48852 36966
rect 21174 36864 21180 36916
rect 21232 36904 21238 36916
rect 24213 36907 24271 36913
rect 24213 36904 24225 36907
rect 21232 36876 24225 36904
rect 21232 36864 21238 36876
rect 24213 36873 24225 36876
rect 24259 36873 24271 36907
rect 25774 36904 25780 36916
rect 25735 36876 25780 36904
rect 24213 36867 24271 36873
rect 25774 36864 25780 36876
rect 25832 36864 25838 36916
rect 29362 36864 29368 36916
rect 29420 36904 29426 36916
rect 29641 36907 29699 36913
rect 29641 36904 29653 36907
rect 29420 36876 29653 36904
rect 29420 36864 29426 36876
rect 29641 36873 29653 36876
rect 29687 36873 29699 36907
rect 47670 36904 47676 36916
rect 47631 36876 47676 36904
rect 29641 36867 29699 36873
rect 47670 36864 47676 36876
rect 47728 36864 47734 36916
rect 7374 36836 7380 36848
rect 7335 36808 7380 36836
rect 7374 36796 7380 36808
rect 7432 36796 7438 36848
rect 17402 36796 17408 36848
rect 17460 36836 17466 36848
rect 20533 36839 20591 36845
rect 20533 36836 20545 36839
rect 17460 36808 20545 36836
rect 17460 36796 17466 36808
rect 20533 36805 20545 36808
rect 20579 36805 20591 36839
rect 20533 36799 20591 36805
rect 23845 36839 23903 36845
rect 23845 36805 23857 36839
rect 23891 36836 23903 36839
rect 24394 36836 24400 36848
rect 23891 36808 24400 36836
rect 23891 36805 23903 36808
rect 23845 36799 23903 36805
rect 24394 36796 24400 36808
rect 24452 36796 24458 36848
rect 24578 36796 24584 36848
rect 24636 36836 24642 36848
rect 46382 36836 46388 36848
rect 24636 36808 46388 36836
rect 24636 36796 24642 36808
rect 46382 36796 46388 36808
rect 46440 36836 46446 36848
rect 46440 36808 47624 36836
rect 46440 36796 46446 36808
rect 18046 36768 18052 36780
rect 18007 36740 18052 36768
rect 18046 36728 18052 36740
rect 18104 36728 18110 36780
rect 18141 36771 18199 36777
rect 18141 36737 18153 36771
rect 18187 36737 18199 36771
rect 18141 36731 18199 36737
rect 7193 36703 7251 36709
rect 7193 36669 7205 36703
rect 7239 36700 7251 36703
rect 8202 36700 8208 36712
rect 7239 36672 8208 36700
rect 7239 36669 7251 36672
rect 7193 36663 7251 36669
rect 8202 36660 8208 36672
rect 8260 36660 8266 36712
rect 8294 36660 8300 36712
rect 8352 36700 8358 36712
rect 8352 36672 8397 36700
rect 8352 36660 8358 36672
rect 17126 36592 17132 36644
rect 17184 36632 17190 36644
rect 18046 36632 18052 36644
rect 17184 36604 18052 36632
rect 17184 36592 17190 36604
rect 18046 36592 18052 36604
rect 18104 36632 18110 36644
rect 18156 36632 18184 36731
rect 18230 36728 18236 36780
rect 18288 36768 18294 36780
rect 18417 36771 18475 36777
rect 18288 36740 18333 36768
rect 18288 36728 18294 36740
rect 18417 36737 18429 36771
rect 18463 36737 18475 36771
rect 18417 36731 18475 36737
rect 18322 36660 18328 36712
rect 18380 36700 18386 36712
rect 18432 36700 18460 36731
rect 19334 36728 19340 36780
rect 19392 36768 19398 36780
rect 19613 36771 19671 36777
rect 19613 36768 19625 36771
rect 19392 36740 19625 36768
rect 19392 36728 19398 36740
rect 19613 36737 19625 36740
rect 19659 36737 19671 36771
rect 19613 36731 19671 36737
rect 19705 36771 19763 36777
rect 19705 36737 19717 36771
rect 19751 36768 19763 36771
rect 23566 36768 23572 36780
rect 19751 36740 23572 36768
rect 19751 36737 19763 36740
rect 19705 36731 19763 36737
rect 23566 36728 23572 36740
rect 23624 36728 23630 36780
rect 23750 36728 23756 36780
rect 23808 36768 23814 36780
rect 24029 36771 24087 36777
rect 24029 36768 24041 36771
rect 23808 36740 24041 36768
rect 23808 36728 23814 36740
rect 24029 36737 24041 36740
rect 24075 36737 24087 36771
rect 24029 36731 24087 36737
rect 25685 36771 25743 36777
rect 25685 36737 25697 36771
rect 25731 36768 25743 36771
rect 25866 36768 25872 36780
rect 25731 36740 25872 36768
rect 25731 36737 25743 36740
rect 25685 36731 25743 36737
rect 25866 36728 25872 36740
rect 25924 36728 25930 36780
rect 26970 36728 26976 36780
rect 27028 36768 27034 36780
rect 27065 36771 27123 36777
rect 27065 36768 27077 36771
rect 27028 36740 27077 36768
rect 27028 36728 27034 36740
rect 27065 36737 27077 36740
rect 27111 36737 27123 36771
rect 27798 36768 27804 36780
rect 27759 36740 27804 36768
rect 27065 36731 27123 36737
rect 27798 36728 27804 36740
rect 27856 36728 27862 36780
rect 27890 36728 27896 36780
rect 27948 36768 27954 36780
rect 28057 36771 28115 36777
rect 28057 36768 28069 36771
rect 27948 36740 28069 36768
rect 27948 36728 27954 36740
rect 28057 36737 28069 36740
rect 28103 36737 28115 36771
rect 29822 36768 29828 36780
rect 29783 36740 29828 36768
rect 28057 36731 28115 36737
rect 29822 36728 29828 36740
rect 29880 36728 29886 36780
rect 30006 36768 30012 36780
rect 29967 36740 30012 36768
rect 30006 36728 30012 36740
rect 30064 36728 30070 36780
rect 30101 36771 30159 36777
rect 30101 36737 30113 36771
rect 30147 36768 30159 36771
rect 30926 36768 30932 36780
rect 30147 36740 30932 36768
rect 30147 36737 30159 36740
rect 30101 36731 30159 36737
rect 19886 36700 19892 36712
rect 18380 36672 18460 36700
rect 19847 36672 19892 36700
rect 18380 36660 18386 36672
rect 19886 36660 19892 36672
rect 19944 36660 19950 36712
rect 20990 36700 20996 36712
rect 19987 36672 20996 36700
rect 19987 36632 20015 36672
rect 20990 36660 20996 36672
rect 21048 36660 21054 36712
rect 25961 36703 26019 36709
rect 25961 36669 25973 36703
rect 26007 36700 26019 36703
rect 26142 36700 26148 36712
rect 26007 36672 26148 36700
rect 26007 36669 26019 36672
rect 25961 36663 26019 36669
rect 26142 36660 26148 36672
rect 26200 36660 26206 36712
rect 30116 36700 30144 36731
rect 30926 36728 30932 36740
rect 30984 36728 30990 36780
rect 46290 36728 46296 36780
rect 46348 36768 46354 36780
rect 47596 36777 47624 36808
rect 47029 36771 47087 36777
rect 47029 36768 47041 36771
rect 46348 36740 47041 36768
rect 46348 36728 46354 36740
rect 47029 36737 47041 36740
rect 47075 36737 47087 36771
rect 47029 36731 47087 36737
rect 47581 36771 47639 36777
rect 47581 36737 47593 36771
rect 47627 36737 47639 36771
rect 47581 36731 47639 36737
rect 29104 36672 30144 36700
rect 18104 36604 20015 36632
rect 18104 36592 18110 36604
rect 20622 36592 20628 36644
rect 20680 36632 20686 36644
rect 20717 36635 20775 36641
rect 20717 36632 20729 36635
rect 20680 36604 20729 36632
rect 20680 36592 20686 36604
rect 20717 36601 20729 36604
rect 20763 36601 20775 36635
rect 20717 36595 20775 36601
rect 23566 36592 23572 36644
rect 23624 36632 23630 36644
rect 23624 36604 27292 36632
rect 23624 36592 23630 36604
rect 2038 36524 2044 36576
rect 2096 36564 2102 36576
rect 2317 36567 2375 36573
rect 2317 36564 2329 36567
rect 2096 36536 2329 36564
rect 2096 36524 2102 36536
rect 2317 36533 2329 36536
rect 2363 36533 2375 36567
rect 2317 36527 2375 36533
rect 17773 36567 17831 36573
rect 17773 36533 17785 36567
rect 17819 36564 17831 36567
rect 18138 36564 18144 36576
rect 17819 36536 18144 36564
rect 17819 36533 17831 36536
rect 17773 36527 17831 36533
rect 18138 36524 18144 36536
rect 18196 36524 18202 36576
rect 19242 36564 19248 36576
rect 19203 36536 19248 36564
rect 19242 36524 19248 36536
rect 19300 36524 19306 36576
rect 20898 36524 20904 36576
rect 20956 36564 20962 36576
rect 24578 36564 24584 36576
rect 20956 36536 24584 36564
rect 20956 36524 20962 36536
rect 24578 36524 24584 36536
rect 24636 36524 24642 36576
rect 25317 36567 25375 36573
rect 25317 36533 25329 36567
rect 25363 36564 25375 36567
rect 25958 36564 25964 36576
rect 25363 36536 25964 36564
rect 25363 36533 25375 36536
rect 25317 36527 25375 36533
rect 25958 36524 25964 36536
rect 26016 36524 26022 36576
rect 26326 36524 26332 36576
rect 26384 36564 26390 36576
rect 27062 36564 27068 36576
rect 26384 36536 27068 36564
rect 26384 36524 26390 36536
rect 27062 36524 27068 36536
rect 27120 36564 27126 36576
rect 27157 36567 27215 36573
rect 27157 36564 27169 36567
rect 27120 36536 27169 36564
rect 27120 36524 27126 36536
rect 27157 36533 27169 36536
rect 27203 36533 27215 36567
rect 27264 36564 27292 36604
rect 29104 36564 29132 36672
rect 27264 36536 29132 36564
rect 29181 36567 29239 36573
rect 27157 36527 27215 36533
rect 29181 36533 29193 36567
rect 29227 36564 29239 36567
rect 29638 36564 29644 36576
rect 29227 36536 29644 36564
rect 29227 36533 29239 36536
rect 29181 36527 29239 36533
rect 29638 36524 29644 36536
rect 29696 36524 29702 36576
rect 1104 36474 48852 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 48852 36474
rect 1104 36400 48852 36422
rect 3326 36320 3332 36372
rect 3384 36360 3390 36372
rect 8202 36360 8208 36372
rect 3384 36332 7788 36360
rect 8163 36332 8208 36360
rect 3384 36320 3390 36332
rect 7760 36292 7788 36332
rect 8202 36320 8208 36332
rect 8260 36320 8266 36372
rect 17126 36360 17132 36372
rect 17087 36332 17132 36360
rect 17126 36320 17132 36332
rect 17184 36320 17190 36372
rect 17678 36360 17684 36372
rect 17639 36332 17684 36360
rect 17678 36320 17684 36332
rect 17736 36320 17742 36372
rect 18230 36320 18236 36372
rect 18288 36360 18294 36372
rect 19613 36363 19671 36369
rect 19613 36360 19625 36363
rect 18288 36332 19625 36360
rect 18288 36320 18294 36332
rect 19613 36329 19625 36332
rect 19659 36329 19671 36363
rect 19613 36323 19671 36329
rect 19886 36320 19892 36372
rect 19944 36360 19950 36372
rect 19944 36332 22094 36360
rect 19944 36320 19950 36332
rect 7760 36264 19334 36292
rect 18598 36224 18604 36236
rect 18156 36196 18604 36224
rect 2961 36159 3019 36165
rect 2961 36125 2973 36159
rect 3007 36156 3019 36159
rect 3326 36156 3332 36168
rect 3007 36128 3332 36156
rect 3007 36125 3019 36128
rect 2961 36119 3019 36125
rect 3326 36116 3332 36128
rect 3384 36116 3390 36168
rect 6825 36159 6883 36165
rect 6825 36125 6837 36159
rect 6871 36156 6883 36159
rect 15562 36156 15568 36168
rect 6871 36128 15568 36156
rect 6871 36125 6883 36128
rect 6825 36119 6883 36125
rect 15562 36116 15568 36128
rect 15620 36116 15626 36168
rect 17034 36156 17040 36168
rect 16995 36128 17040 36156
rect 17034 36116 17040 36128
rect 17092 36116 17098 36168
rect 17678 36116 17684 36168
rect 17736 36156 17742 36168
rect 18156 36165 18184 36196
rect 18598 36184 18604 36196
rect 18656 36184 18662 36236
rect 19306 36224 19334 36264
rect 20070 36252 20076 36304
rect 20128 36292 20134 36304
rect 20438 36292 20444 36304
rect 20128 36264 20444 36292
rect 20128 36252 20134 36264
rect 20438 36252 20444 36264
rect 20496 36252 20502 36304
rect 21637 36295 21695 36301
rect 21637 36261 21649 36295
rect 21683 36261 21695 36295
rect 21637 36255 21695 36261
rect 20898 36224 20904 36236
rect 19306 36196 20904 36224
rect 17911 36159 17969 36165
rect 17911 36156 17923 36159
rect 17736 36128 17923 36156
rect 17736 36116 17742 36128
rect 17911 36125 17923 36128
rect 17957 36125 17969 36159
rect 17911 36119 17969 36125
rect 18046 36156 18104 36162
rect 18046 36122 18058 36156
rect 18092 36122 18104 36156
rect 18046 36116 18104 36122
rect 18141 36159 18199 36165
rect 18141 36125 18153 36159
rect 18187 36125 18199 36159
rect 18322 36156 18328 36168
rect 18283 36128 18328 36156
rect 18141 36119 18199 36125
rect 18322 36116 18328 36128
rect 18380 36116 18386 36168
rect 19242 36156 19248 36168
rect 19203 36128 19248 36156
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 19426 36156 19432 36168
rect 19387 36128 19432 36156
rect 19426 36116 19432 36128
rect 19484 36116 19490 36168
rect 20180 36165 20208 36196
rect 20898 36184 20904 36196
rect 20956 36184 20962 36236
rect 20165 36159 20223 36165
rect 20165 36125 20177 36159
rect 20211 36125 20223 36159
rect 20165 36119 20223 36125
rect 20809 36159 20867 36165
rect 20809 36125 20821 36159
rect 20855 36156 20867 36159
rect 21652 36156 21680 36255
rect 22066 36224 22094 36332
rect 22186 36320 22192 36372
rect 22244 36360 22250 36372
rect 24857 36363 24915 36369
rect 24857 36360 24869 36363
rect 22244 36332 24869 36360
rect 22244 36320 22250 36332
rect 24857 36329 24869 36332
rect 24903 36329 24915 36363
rect 24857 36323 24915 36329
rect 26881 36363 26939 36369
rect 26881 36329 26893 36363
rect 26927 36360 26939 36363
rect 27890 36360 27896 36372
rect 26927 36332 27896 36360
rect 26927 36329 26939 36332
rect 26881 36323 26939 36329
rect 27890 36320 27896 36332
rect 27948 36320 27954 36372
rect 22462 36252 22468 36304
rect 22520 36292 22526 36304
rect 26786 36292 26792 36304
rect 22520 36264 26792 36292
rect 22520 36252 22526 36264
rect 26786 36252 26792 36264
rect 26844 36292 26850 36304
rect 26844 36264 27261 36292
rect 26844 36252 26850 36264
rect 22281 36227 22339 36233
rect 22281 36224 22293 36227
rect 22066 36196 22293 36224
rect 22281 36193 22293 36196
rect 22327 36224 22339 36227
rect 22327 36196 23244 36224
rect 22327 36193 22339 36196
rect 22281 36187 22339 36193
rect 20855 36128 21680 36156
rect 22097 36159 22155 36165
rect 20855 36125 20867 36128
rect 20809 36119 20867 36125
rect 22097 36125 22109 36159
rect 22143 36156 22155 36159
rect 23106 36156 23112 36168
rect 22143 36128 23112 36156
rect 22143 36125 22155 36128
rect 22097 36119 22155 36125
rect 23106 36116 23112 36128
rect 23164 36116 23170 36168
rect 7092 36091 7150 36097
rect 7092 36057 7104 36091
rect 7138 36088 7150 36091
rect 7650 36088 7656 36100
rect 7138 36060 7656 36088
rect 7138 36057 7150 36060
rect 7092 36051 7150 36057
rect 7650 36048 7656 36060
rect 7708 36048 7714 36100
rect 3050 36020 3056 36032
rect 3011 35992 3056 36020
rect 3050 35980 3056 35992
rect 3108 35980 3114 36032
rect 18064 36020 18092 36116
rect 19444 36088 19472 36116
rect 20993 36091 21051 36097
rect 20993 36088 21005 36091
rect 19444 36060 21005 36088
rect 20993 36057 21005 36060
rect 21039 36057 21051 36091
rect 20993 36051 21051 36057
rect 23216 36032 23244 36196
rect 24765 36159 24823 36165
rect 24765 36125 24777 36159
rect 24811 36156 24823 36159
rect 26326 36156 26332 36168
rect 24811 36128 26332 36156
rect 24811 36125 24823 36128
rect 24765 36119 24823 36125
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 27233 36165 27261 36264
rect 28166 36252 28172 36304
rect 28224 36292 28230 36304
rect 30006 36292 30012 36304
rect 28224 36264 30012 36292
rect 28224 36252 28230 36264
rect 30006 36252 30012 36264
rect 30064 36252 30070 36304
rect 27137 36159 27195 36165
rect 27137 36125 27149 36159
rect 27183 36156 27195 36159
rect 27230 36159 27288 36165
rect 27183 36125 27200 36156
rect 27137 36119 27200 36125
rect 27230 36125 27242 36159
rect 27276 36125 27288 36159
rect 27230 36119 27288 36125
rect 27341 36156 27399 36162
rect 27522 36156 27528 36168
rect 27341 36122 27353 36156
rect 27387 36122 27399 36156
rect 27483 36128 27528 36156
rect 23569 36091 23627 36097
rect 23569 36057 23581 36091
rect 23615 36088 23627 36091
rect 24394 36088 24400 36100
rect 23615 36060 24400 36088
rect 23615 36057 23627 36060
rect 23569 36051 23627 36057
rect 24394 36048 24400 36060
rect 24452 36048 24458 36100
rect 25958 36088 25964 36100
rect 25919 36060 25964 36088
rect 25958 36048 25964 36060
rect 26016 36048 26022 36100
rect 26145 36091 26203 36097
rect 26145 36057 26157 36091
rect 26191 36057 26203 36091
rect 26145 36051 26203 36057
rect 18506 36020 18512 36032
rect 18064 35992 18512 36020
rect 18506 35980 18512 35992
rect 18564 35980 18570 36032
rect 20070 35980 20076 36032
rect 20128 36020 20134 36032
rect 20257 36023 20315 36029
rect 20257 36020 20269 36023
rect 20128 35992 20269 36020
rect 20128 35980 20134 35992
rect 20257 35989 20269 35992
rect 20303 35989 20315 36023
rect 20257 35983 20315 35989
rect 21082 35980 21088 36032
rect 21140 36020 21146 36032
rect 21177 36023 21235 36029
rect 21177 36020 21189 36023
rect 21140 35992 21189 36020
rect 21140 35980 21146 35992
rect 21177 35989 21189 35992
rect 21223 35989 21235 36023
rect 21177 35983 21235 35989
rect 22005 36023 22063 36029
rect 22005 35989 22017 36023
rect 22051 36020 22063 36023
rect 23106 36020 23112 36032
rect 22051 35992 23112 36020
rect 22051 35989 22063 35992
rect 22005 35983 22063 35989
rect 23106 35980 23112 35992
rect 23164 35980 23170 36032
rect 23198 35980 23204 36032
rect 23256 36020 23262 36032
rect 23661 36023 23719 36029
rect 23661 36020 23673 36023
rect 23256 35992 23673 36020
rect 23256 35980 23262 35992
rect 23661 35989 23673 35992
rect 23707 35989 23719 36023
rect 23661 35983 23719 35989
rect 24578 35980 24584 36032
rect 24636 36020 24642 36032
rect 26160 36020 26188 36051
rect 26878 36048 26884 36100
rect 26936 36088 26942 36100
rect 27172 36088 27200 36119
rect 27341 36116 27399 36122
rect 27522 36116 27528 36128
rect 27580 36116 27586 36168
rect 47854 36156 47860 36168
rect 47815 36128 47860 36156
rect 47854 36116 47860 36128
rect 47912 36116 47918 36168
rect 26936 36060 27200 36088
rect 26936 36048 26942 36060
rect 24636 35992 26188 36020
rect 26329 36023 26387 36029
rect 24636 35980 24642 35992
rect 26329 35989 26341 36023
rect 26375 36020 26387 36023
rect 27356 36020 27384 36116
rect 26375 35992 27384 36020
rect 48041 36023 48099 36029
rect 26375 35989 26387 35992
rect 26329 35983 26387 35989
rect 48041 35989 48053 36023
rect 48087 36020 48099 36023
rect 48130 36020 48136 36032
rect 48087 35992 48136 36020
rect 48087 35989 48099 35992
rect 48041 35983 48099 35989
rect 48130 35980 48136 35992
rect 48188 35980 48194 36032
rect 1104 35930 48852 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 48852 35930
rect 1104 35856 48852 35878
rect 1578 35776 1584 35828
rect 1636 35816 1642 35828
rect 7650 35816 7656 35828
rect 1636 35788 7512 35816
rect 7611 35788 7656 35816
rect 1636 35776 1642 35788
rect 2225 35751 2283 35757
rect 2225 35717 2237 35751
rect 2271 35748 2283 35751
rect 3050 35748 3056 35760
rect 2271 35720 3056 35748
rect 2271 35717 2283 35720
rect 2225 35711 2283 35717
rect 3050 35708 3056 35720
rect 3108 35708 3114 35760
rect 7484 35748 7512 35788
rect 7650 35776 7656 35788
rect 7708 35776 7714 35828
rect 8386 35776 8392 35828
rect 8444 35816 8450 35828
rect 24670 35816 24676 35828
rect 8444 35788 24676 35816
rect 8444 35776 8450 35788
rect 24670 35776 24676 35788
rect 24728 35776 24734 35828
rect 25593 35819 25651 35825
rect 25593 35816 25605 35819
rect 24780 35788 25605 35816
rect 17402 35748 17408 35760
rect 7484 35720 12434 35748
rect 17363 35720 17408 35748
rect 2038 35680 2044 35692
rect 1999 35652 2044 35680
rect 2038 35640 2044 35652
rect 2096 35640 2102 35692
rect 7837 35683 7895 35689
rect 7837 35649 7849 35683
rect 7883 35649 7895 35683
rect 7837 35643 7895 35649
rect 2774 35572 2780 35624
rect 2832 35612 2838 35624
rect 2832 35584 2877 35612
rect 2832 35572 2838 35584
rect 7852 35476 7880 35643
rect 12406 35544 12434 35720
rect 17402 35708 17408 35720
rect 17460 35708 17466 35760
rect 18322 35708 18328 35760
rect 18380 35748 18386 35760
rect 19886 35748 19892 35760
rect 18380 35720 19892 35748
rect 18380 35708 18386 35720
rect 19886 35708 19892 35720
rect 19944 35708 19950 35760
rect 20625 35751 20683 35757
rect 20625 35717 20637 35751
rect 20671 35748 20683 35751
rect 20714 35748 20720 35760
rect 20671 35720 20720 35748
rect 20671 35717 20683 35720
rect 20625 35711 20683 35717
rect 20714 35708 20720 35720
rect 20772 35708 20778 35760
rect 22186 35748 22192 35760
rect 21836 35720 22192 35748
rect 17221 35683 17279 35689
rect 17221 35649 17233 35683
rect 17267 35680 17279 35683
rect 17954 35680 17960 35692
rect 17267 35652 17960 35680
rect 17267 35649 17279 35652
rect 17221 35643 17279 35649
rect 17954 35640 17960 35652
rect 18012 35640 18018 35692
rect 18138 35689 18144 35692
rect 18132 35680 18144 35689
rect 18099 35652 18144 35680
rect 18132 35643 18144 35652
rect 18138 35640 18144 35643
rect 18196 35640 18202 35692
rect 20806 35640 20812 35692
rect 20864 35689 20870 35692
rect 20990 35689 20996 35692
rect 20864 35683 20913 35689
rect 20864 35649 20867 35683
rect 20901 35649 20913 35683
rect 20864 35643 20913 35649
rect 20974 35683 20996 35689
rect 20974 35649 20986 35683
rect 20974 35643 20996 35649
rect 20864 35640 20870 35643
rect 20990 35640 20996 35643
rect 21048 35640 21054 35692
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 21269 35686 21327 35689
rect 21269 35683 21404 35686
rect 21140 35652 21185 35680
rect 21140 35640 21146 35652
rect 21269 35649 21281 35683
rect 21315 35680 21404 35683
rect 21450 35680 21456 35692
rect 21315 35658 21456 35680
rect 21315 35649 21327 35658
rect 21376 35652 21456 35658
rect 21269 35643 21327 35649
rect 21450 35640 21456 35652
rect 21508 35640 21514 35692
rect 21836 35689 21864 35720
rect 22186 35708 22192 35720
rect 22244 35708 22250 35760
rect 24121 35751 24179 35757
rect 24121 35717 24133 35751
rect 24167 35748 24179 35751
rect 24210 35748 24216 35760
rect 24167 35720 24216 35748
rect 24167 35717 24179 35720
rect 24121 35711 24179 35717
rect 24210 35708 24216 35720
rect 24268 35708 24274 35760
rect 24780 35757 24808 35788
rect 25593 35785 25605 35788
rect 25639 35785 25651 35819
rect 25593 35779 25651 35785
rect 25774 35776 25780 35828
rect 25832 35816 25838 35828
rect 25961 35819 26019 35825
rect 25961 35816 25973 35819
rect 25832 35788 25973 35816
rect 25832 35776 25838 35788
rect 25961 35785 25973 35788
rect 26007 35816 26019 35819
rect 28721 35819 28779 35825
rect 28721 35816 28733 35819
rect 26007 35788 28733 35816
rect 26007 35785 26019 35788
rect 25961 35779 26019 35785
rect 28721 35785 28733 35788
rect 28767 35785 28779 35819
rect 28721 35779 28779 35785
rect 24765 35751 24823 35757
rect 24765 35717 24777 35751
rect 24811 35717 24823 35751
rect 26053 35751 26111 35757
rect 26053 35748 26065 35751
rect 24765 35711 24823 35717
rect 24872 35720 26065 35748
rect 21821 35683 21879 35689
rect 21821 35649 21833 35683
rect 21867 35649 21879 35683
rect 21821 35643 21879 35649
rect 21910 35640 21916 35692
rect 21968 35680 21974 35692
rect 22077 35683 22135 35689
rect 22077 35680 22089 35683
rect 21968 35652 22089 35680
rect 21968 35640 21974 35652
rect 22077 35649 22089 35652
rect 22123 35649 22135 35683
rect 22077 35643 22135 35649
rect 23658 35640 23664 35692
rect 23716 35680 23722 35692
rect 23937 35683 23995 35689
rect 23937 35680 23949 35683
rect 23716 35652 23949 35680
rect 23716 35640 23722 35652
rect 23937 35649 23949 35652
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 24486 35640 24492 35692
rect 24544 35680 24550 35692
rect 24872 35680 24900 35720
rect 26053 35717 26065 35720
rect 26099 35717 26111 35751
rect 27798 35748 27804 35760
rect 26053 35711 26111 35717
rect 27356 35720 27804 35748
rect 27356 35689 27384 35720
rect 27798 35708 27804 35720
rect 27856 35708 27862 35760
rect 24544 35652 24900 35680
rect 24949 35683 25007 35689
rect 24544 35640 24550 35652
rect 24949 35649 24961 35683
rect 24995 35649 25007 35683
rect 24949 35643 25007 35649
rect 27341 35683 27399 35689
rect 27341 35649 27353 35683
rect 27387 35649 27399 35683
rect 27341 35643 27399 35649
rect 15562 35572 15568 35624
rect 15620 35612 15626 35624
rect 16482 35612 16488 35624
rect 15620 35584 16488 35612
rect 15620 35572 15626 35584
rect 16482 35572 16488 35584
rect 16540 35612 16546 35624
rect 17865 35615 17923 35621
rect 17865 35612 17877 35615
rect 16540 35584 17877 35612
rect 16540 35572 16546 35584
rect 17865 35581 17877 35584
rect 17911 35581 17923 35615
rect 17865 35575 17923 35581
rect 23750 35572 23756 35624
rect 23808 35612 23814 35624
rect 24578 35612 24584 35624
rect 23808 35584 24584 35612
rect 23808 35572 23814 35584
rect 24578 35572 24584 35584
rect 24636 35612 24642 35624
rect 24964 35612 24992 35643
rect 27430 35640 27436 35692
rect 27488 35680 27494 35692
rect 27597 35683 27655 35689
rect 27597 35680 27609 35683
rect 27488 35652 27609 35680
rect 27488 35640 27494 35652
rect 27597 35649 27609 35652
rect 27643 35649 27655 35683
rect 27597 35643 27655 35649
rect 48222 35640 48228 35692
rect 48280 35640 48286 35692
rect 26234 35612 26240 35624
rect 24636 35584 24992 35612
rect 26195 35584 26240 35612
rect 24636 35572 24642 35584
rect 26234 35572 26240 35584
rect 26292 35572 26298 35624
rect 27338 35544 27344 35556
rect 12406 35516 17264 35544
rect 17126 35476 17132 35488
rect 7852 35448 17132 35476
rect 17126 35436 17132 35448
rect 17184 35436 17190 35488
rect 17236 35476 17264 35516
rect 18800 35516 20760 35544
rect 18800 35476 18828 35516
rect 17236 35448 18828 35476
rect 19245 35479 19303 35485
rect 19245 35445 19257 35479
rect 19291 35476 19303 35479
rect 19334 35476 19340 35488
rect 19291 35448 19340 35476
rect 19291 35445 19303 35448
rect 19245 35439 19303 35445
rect 19334 35436 19340 35448
rect 19392 35476 19398 35488
rect 19794 35476 19800 35488
rect 19392 35448 19800 35476
rect 19392 35436 19398 35448
rect 19794 35436 19800 35448
rect 19852 35436 19858 35488
rect 20732 35476 20760 35516
rect 23124 35516 27344 35544
rect 23124 35476 23152 35516
rect 27338 35504 27344 35516
rect 27396 35504 27402 35556
rect 48240 35488 48268 35640
rect 20732 35448 23152 35476
rect 23201 35479 23259 35485
rect 23201 35445 23213 35479
rect 23247 35476 23259 35479
rect 23290 35476 23296 35488
rect 23247 35448 23296 35476
rect 23247 35445 23259 35448
rect 23201 35439 23259 35445
rect 23290 35436 23296 35448
rect 23348 35436 23354 35488
rect 25133 35479 25191 35485
rect 25133 35445 25145 35479
rect 25179 35476 25191 35479
rect 27246 35476 27252 35488
rect 25179 35448 27252 35476
rect 25179 35445 25191 35448
rect 25133 35439 25191 35445
rect 27246 35436 27252 35448
rect 27304 35436 27310 35488
rect 47210 35436 47216 35488
rect 47268 35476 47274 35488
rect 47765 35479 47823 35485
rect 47765 35476 47777 35479
rect 47268 35448 47777 35476
rect 47268 35436 47274 35448
rect 47765 35445 47777 35448
rect 47811 35445 47823 35479
rect 47765 35439 47823 35445
rect 48222 35436 48228 35488
rect 48280 35436 48286 35488
rect 1104 35386 48852 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 48852 35386
rect 1104 35312 48852 35334
rect 15562 35272 15568 35284
rect 15523 35244 15568 35272
rect 15562 35232 15568 35244
rect 15620 35232 15626 35284
rect 24578 35272 24584 35284
rect 20548 35244 22048 35272
rect 24539 35244 24584 35272
rect 2746 35176 17540 35204
rect 1673 35139 1731 35145
rect 1673 35105 1685 35139
rect 1719 35136 1731 35139
rect 2746 35136 2774 35176
rect 1719 35108 2774 35136
rect 11425 35139 11483 35145
rect 1719 35105 1731 35108
rect 1673 35099 1731 35105
rect 11425 35105 11437 35139
rect 11471 35136 11483 35139
rect 13078 35136 13084 35148
rect 11471 35108 13084 35136
rect 11471 35105 11483 35108
rect 11425 35099 11483 35105
rect 13078 35096 13084 35108
rect 13136 35096 13142 35148
rect 13262 35136 13268 35148
rect 13223 35108 13268 35136
rect 13262 35096 13268 35108
rect 13320 35096 13326 35148
rect 1394 35068 1400 35080
rect 1355 35040 1400 35068
rect 1394 35028 1400 35040
rect 1452 35028 1458 35080
rect 15473 35071 15531 35077
rect 15473 35037 15485 35071
rect 15519 35068 15531 35071
rect 17402 35068 17408 35080
rect 15519 35040 17408 35068
rect 15519 35037 15531 35040
rect 15473 35031 15531 35037
rect 17402 35028 17408 35040
rect 17460 35028 17466 35080
rect 17512 35068 17540 35176
rect 17678 35164 17684 35216
rect 17736 35204 17742 35216
rect 18966 35204 18972 35216
rect 17736 35176 18972 35204
rect 17736 35164 17742 35176
rect 18966 35164 18972 35176
rect 19024 35164 19030 35216
rect 19889 35139 19947 35145
rect 19889 35105 19901 35139
rect 19935 35136 19947 35139
rect 19978 35136 19984 35148
rect 19935 35108 19984 35136
rect 19935 35105 19947 35108
rect 19889 35099 19947 35105
rect 19978 35096 19984 35108
rect 20036 35096 20042 35148
rect 20548 35136 20576 35244
rect 20809 35207 20867 35213
rect 20809 35173 20821 35207
rect 20855 35204 20867 35207
rect 22020 35204 22048 35244
rect 24578 35232 24584 35244
rect 24636 35232 24642 35284
rect 26789 35275 26847 35281
rect 26789 35241 26801 35275
rect 26835 35272 26847 35275
rect 27430 35272 27436 35284
rect 26835 35244 27436 35272
rect 26835 35241 26847 35244
rect 26789 35235 26847 35241
rect 27430 35232 27436 35244
rect 27488 35232 27494 35284
rect 27614 35232 27620 35284
rect 27672 35272 27678 35284
rect 28077 35275 28135 35281
rect 28077 35272 28089 35275
rect 27672 35244 28089 35272
rect 27672 35232 27678 35244
rect 28077 35241 28089 35244
rect 28123 35241 28135 35275
rect 28077 35235 28135 35241
rect 22557 35207 22615 35213
rect 22557 35204 22569 35207
rect 20855 35176 21772 35204
rect 22020 35176 22569 35204
rect 20855 35173 20867 35176
rect 20809 35167 20867 35173
rect 21266 35136 21272 35148
rect 20456 35108 20576 35136
rect 21008 35108 21272 35136
rect 17911 35071 17969 35077
rect 17911 35068 17923 35071
rect 17512 35040 17923 35068
rect 17911 35037 17923 35040
rect 17957 35037 17969 35071
rect 18043 35068 18049 35080
rect 18004 35040 18049 35068
rect 17911 35031 17969 35037
rect 18043 35028 18049 35040
rect 18101 35028 18107 35080
rect 18138 35028 18144 35080
rect 18196 35077 18202 35080
rect 18196 35068 18204 35077
rect 18322 35068 18328 35080
rect 18196 35040 18241 35068
rect 18283 35040 18328 35068
rect 18196 35031 18204 35040
rect 18196 35028 18202 35031
rect 18322 35028 18328 35040
rect 18380 35028 18386 35080
rect 19334 35028 19340 35080
rect 19392 35068 19398 35080
rect 19610 35068 19616 35080
rect 19392 35040 19616 35068
rect 19392 35028 19398 35040
rect 19610 35028 19616 35040
rect 19668 35028 19674 35080
rect 20456 35077 20484 35108
rect 20441 35071 20499 35077
rect 20441 35037 20453 35071
rect 20487 35037 20499 35071
rect 21008 35068 21036 35108
rect 21266 35096 21272 35108
rect 21324 35096 21330 35148
rect 21542 35077 21548 35080
rect 20441 35031 20499 35037
rect 20548 35040 21036 35068
rect 21525 35071 21548 35077
rect 11606 35000 11612 35012
rect 11567 34972 11612 35000
rect 11606 34960 11612 34972
rect 11664 34960 11670 35012
rect 19705 35003 19763 35009
rect 19705 34969 19717 35003
rect 19751 35000 19763 35003
rect 20548 35000 20576 35040
rect 21525 35037 21537 35071
rect 21525 35031 21548 35037
rect 21542 35028 21548 35031
rect 21600 35028 21606 35080
rect 21744 35077 21772 35176
rect 22557 35173 22569 35176
rect 22603 35173 22615 35207
rect 22557 35167 22615 35173
rect 24670 35164 24676 35216
rect 24728 35204 24734 35216
rect 24728 35176 31754 35204
rect 24728 35164 24734 35176
rect 23198 35136 23204 35148
rect 23159 35108 23204 35136
rect 23198 35096 23204 35108
rect 23256 35096 23262 35148
rect 23290 35096 23296 35148
rect 23348 35136 23354 35148
rect 24489 35139 24547 35145
rect 24489 35136 24501 35139
rect 23348 35108 24501 35136
rect 23348 35096 23354 35108
rect 24489 35105 24501 35108
rect 24535 35105 24547 35139
rect 25498 35136 25504 35148
rect 25459 35108 25504 35136
rect 24489 35099 24547 35105
rect 25498 35096 25504 35108
rect 25556 35096 25562 35148
rect 25682 35136 25688 35148
rect 25643 35108 25688 35136
rect 25682 35096 25688 35108
rect 25740 35096 25746 35148
rect 26786 35096 26792 35148
rect 26844 35136 26850 35148
rect 31726 35136 31754 35176
rect 32769 35139 32827 35145
rect 32769 35136 32781 35139
rect 26844 35108 27200 35136
rect 31726 35108 32781 35136
rect 26844 35096 26850 35108
rect 21637 35071 21695 35077
rect 21637 35037 21649 35071
rect 21683 35037 21695 35071
rect 21637 35031 21695 35037
rect 21729 35071 21787 35077
rect 21729 35037 21741 35071
rect 21775 35037 21787 35071
rect 21910 35068 21916 35080
rect 21871 35040 21916 35068
rect 21729 35031 21787 35037
rect 19751 34972 20576 35000
rect 20625 35003 20683 35009
rect 19751 34969 19763 34972
rect 19705 34963 19763 34969
rect 20625 34969 20637 35003
rect 20671 35000 20683 35003
rect 20714 35000 20720 35012
rect 20671 34972 20720 35000
rect 20671 34969 20683 34972
rect 20625 34963 20683 34969
rect 20714 34960 20720 34972
rect 20772 34960 20778 35012
rect 20990 34960 20996 35012
rect 21048 35000 21054 35012
rect 21652 35000 21680 35031
rect 21910 35028 21916 35040
rect 21968 35028 21974 35080
rect 22002 35028 22008 35080
rect 22060 35068 22066 35080
rect 24673 35071 24731 35077
rect 24673 35068 24685 35071
rect 22060 35040 24685 35068
rect 22060 35028 22066 35040
rect 24673 35037 24685 35040
rect 24719 35037 24731 35071
rect 24673 35031 24731 35037
rect 25593 35071 25651 35077
rect 25593 35037 25605 35071
rect 25639 35068 25651 35071
rect 26234 35068 26240 35080
rect 25639 35040 26240 35068
rect 25639 35037 25651 35040
rect 25593 35031 25651 35037
rect 26234 35028 26240 35040
rect 26292 35028 26298 35080
rect 27172 35077 27200 35108
rect 32769 35105 32781 35108
rect 32815 35105 32827 35139
rect 32769 35099 32827 35105
rect 46293 35139 46351 35145
rect 46293 35105 46305 35139
rect 46339 35136 46351 35139
rect 47026 35136 47032 35148
rect 46339 35108 47032 35136
rect 46339 35105 46351 35108
rect 46293 35099 46351 35105
rect 47026 35096 47032 35108
rect 47084 35096 47090 35148
rect 48130 35136 48136 35148
rect 48091 35108 48136 35136
rect 48130 35096 48136 35108
rect 48188 35096 48194 35148
rect 27065 35071 27123 35077
rect 27065 35037 27077 35071
rect 27111 35037 27123 35071
rect 27065 35031 27123 35037
rect 27154 35071 27212 35077
rect 27154 35037 27166 35071
rect 27200 35037 27212 35071
rect 27154 35031 27212 35037
rect 21048 34972 21680 35000
rect 22925 35003 22983 35009
rect 21048 34960 21054 34972
rect 22925 34969 22937 35003
rect 22971 35000 22983 35003
rect 23474 35000 23480 35012
rect 22971 34972 23480 35000
rect 22971 34969 22983 34972
rect 22925 34963 22983 34969
rect 23474 34960 23480 34972
rect 23532 34960 23538 35012
rect 24397 35003 24455 35009
rect 24397 34969 24409 35003
rect 24443 35000 24455 35003
rect 24486 35000 24492 35012
rect 24443 34972 24492 35000
rect 24443 34969 24455 34972
rect 24397 34963 24455 34969
rect 24486 34960 24492 34972
rect 24544 34960 24550 35012
rect 25130 35000 25136 35012
rect 24780 34972 25136 35000
rect 17678 34932 17684 34944
rect 17639 34904 17684 34932
rect 17678 34892 17684 34904
rect 17736 34892 17742 34944
rect 19242 34932 19248 34944
rect 19203 34904 19248 34932
rect 19242 34892 19248 34904
rect 19300 34892 19306 34944
rect 21269 34935 21327 34941
rect 21269 34901 21281 34935
rect 21315 34932 21327 34935
rect 21910 34932 21916 34944
rect 21315 34904 21916 34932
rect 21315 34901 21327 34904
rect 21269 34895 21327 34901
rect 21910 34892 21916 34904
rect 21968 34892 21974 34944
rect 23017 34935 23075 34941
rect 23017 34901 23029 34935
rect 23063 34932 23075 34935
rect 24780 34932 24808 34972
rect 25130 34960 25136 34972
rect 25188 34960 25194 35012
rect 25317 35003 25375 35009
rect 25317 34969 25329 35003
rect 25363 34969 25375 35003
rect 25317 34963 25375 34969
rect 23063 34904 24808 34932
rect 24857 34935 24915 34941
rect 23063 34901 23075 34904
rect 23017 34895 23075 34901
rect 24857 34901 24869 34935
rect 24903 34932 24915 34935
rect 25332 34932 25360 34963
rect 24903 34904 25360 34932
rect 25409 34935 25467 34941
rect 24903 34901 24915 34904
rect 24857 34895 24915 34901
rect 25409 34901 25421 34935
rect 25455 34932 25467 34935
rect 25590 34932 25596 34944
rect 25455 34904 25596 34932
rect 25455 34901 25467 34904
rect 25409 34895 25467 34901
rect 25590 34892 25596 34904
rect 25648 34892 25654 34944
rect 27080 34932 27108 35031
rect 27246 35028 27252 35080
rect 27304 35068 27310 35080
rect 27433 35071 27491 35077
rect 27304 35040 27349 35068
rect 27304 35028 27310 35040
rect 27433 35037 27445 35071
rect 27479 35068 27491 35071
rect 27522 35068 27528 35080
rect 27479 35040 27528 35068
rect 27479 35037 27491 35040
rect 27433 35031 27491 35037
rect 27522 35028 27528 35040
rect 27580 35028 27586 35080
rect 32306 35068 32312 35080
rect 32267 35040 32312 35068
rect 32306 35028 32312 35040
rect 32364 35028 32370 35080
rect 27982 35000 27988 35012
rect 27943 34972 27988 35000
rect 27982 34960 27988 34972
rect 28040 34960 28046 35012
rect 32493 35003 32551 35009
rect 32493 34969 32505 35003
rect 32539 35000 32551 35003
rect 33410 35000 33416 35012
rect 32539 34972 33416 35000
rect 32539 34969 32551 34972
rect 32493 34963 32551 34969
rect 33410 34960 33416 34972
rect 33468 34960 33474 35012
rect 46474 35000 46480 35012
rect 46435 34972 46480 35000
rect 46474 34960 46480 34972
rect 46532 34960 46538 35012
rect 27522 34932 27528 34944
rect 27080 34904 27528 34932
rect 27522 34892 27528 34904
rect 27580 34892 27586 34944
rect 1104 34842 48852 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 48852 34842
rect 1104 34768 48852 34790
rect 11606 34728 11612 34740
rect 11567 34700 11612 34728
rect 11606 34688 11612 34700
rect 11664 34688 11670 34740
rect 19153 34731 19211 34737
rect 19153 34697 19165 34731
rect 19199 34728 19211 34731
rect 19334 34728 19340 34740
rect 19199 34700 19340 34728
rect 19199 34697 19211 34700
rect 19153 34691 19211 34697
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 19426 34688 19432 34740
rect 19484 34728 19490 34740
rect 19613 34731 19671 34737
rect 19613 34728 19625 34731
rect 19484 34700 19625 34728
rect 19484 34688 19490 34700
rect 19613 34697 19625 34700
rect 19659 34728 19671 34731
rect 20714 34728 20720 34740
rect 19659 34700 20720 34728
rect 19659 34697 19671 34700
rect 19613 34691 19671 34697
rect 20714 34688 20720 34700
rect 20772 34688 20778 34740
rect 22830 34728 22836 34740
rect 21100 34700 22836 34728
rect 17678 34620 17684 34672
rect 17736 34660 17742 34672
rect 21100 34669 21128 34700
rect 22830 34688 22836 34700
rect 22888 34688 22894 34740
rect 23201 34731 23259 34737
rect 23201 34697 23213 34731
rect 23247 34697 23259 34731
rect 23201 34691 23259 34697
rect 18018 34663 18076 34669
rect 18018 34660 18030 34663
rect 17736 34632 18030 34660
rect 17736 34620 17742 34632
rect 18018 34629 18030 34632
rect 18064 34629 18076 34663
rect 18018 34623 18076 34629
rect 21085 34663 21143 34669
rect 21085 34629 21097 34663
rect 21131 34629 21143 34663
rect 22186 34660 22192 34672
rect 21085 34623 21143 34629
rect 21836 34632 22192 34660
rect 11514 34592 11520 34604
rect 11475 34564 11520 34592
rect 11514 34552 11520 34564
rect 11572 34592 11578 34604
rect 11974 34592 11980 34604
rect 11572 34564 11980 34592
rect 11572 34552 11578 34564
rect 11974 34552 11980 34564
rect 12032 34552 12038 34604
rect 15562 34552 15568 34604
rect 15620 34592 15626 34604
rect 17773 34595 17831 34601
rect 17773 34592 17785 34595
rect 15620 34564 17785 34592
rect 15620 34552 15626 34564
rect 17773 34561 17785 34564
rect 17819 34561 17831 34595
rect 17773 34555 17831 34561
rect 19334 34552 19340 34604
rect 19392 34592 19398 34604
rect 21836 34601 21864 34632
rect 22186 34620 22192 34632
rect 22244 34620 22250 34672
rect 23216 34660 23244 34691
rect 24578 34688 24584 34740
rect 24636 34728 24642 34740
rect 25409 34731 25467 34737
rect 25409 34728 25421 34731
rect 24636 34700 25421 34728
rect 24636 34688 24642 34700
rect 25409 34697 25421 34700
rect 25455 34697 25467 34731
rect 25409 34691 25467 34697
rect 26329 34731 26387 34737
rect 26329 34697 26341 34731
rect 26375 34728 26387 34731
rect 26602 34728 26608 34740
rect 26375 34700 26608 34728
rect 26375 34697 26387 34700
rect 26329 34691 26387 34697
rect 26602 34688 26608 34700
rect 26660 34688 26666 34740
rect 32306 34688 32312 34740
rect 32364 34728 32370 34740
rect 33505 34731 33563 34737
rect 33505 34728 33517 34731
rect 32364 34700 33517 34728
rect 32364 34688 32370 34700
rect 33505 34697 33517 34700
rect 33551 34697 33563 34731
rect 33505 34691 33563 34697
rect 23474 34660 23480 34672
rect 23216 34632 23480 34660
rect 23474 34620 23480 34632
rect 23532 34660 23538 34672
rect 24670 34660 24676 34672
rect 23532 34632 24676 34660
rect 23532 34620 23538 34632
rect 24670 34620 24676 34632
rect 24728 34620 24734 34672
rect 26620 34660 26648 34688
rect 26620 34632 27016 34660
rect 19797 34595 19855 34601
rect 19797 34592 19809 34595
rect 19392 34564 19809 34592
rect 19392 34552 19398 34564
rect 19797 34561 19809 34564
rect 19843 34592 19855 34595
rect 21821 34595 21879 34601
rect 19843 34564 21772 34592
rect 19843 34561 19855 34564
rect 19797 34555 19855 34561
rect 21266 34524 21272 34536
rect 21227 34496 21272 34524
rect 21266 34484 21272 34496
rect 21324 34484 21330 34536
rect 21744 34524 21772 34564
rect 21821 34561 21833 34595
rect 21867 34561 21879 34595
rect 21821 34555 21879 34561
rect 21910 34552 21916 34604
rect 21968 34592 21974 34604
rect 22077 34595 22135 34601
rect 22077 34592 22089 34595
rect 21968 34564 22089 34592
rect 21968 34552 21974 34564
rect 22077 34561 22089 34564
rect 22123 34561 22135 34595
rect 25314 34592 25320 34604
rect 25275 34564 25320 34592
rect 22077 34555 22135 34561
rect 25314 34552 25320 34564
rect 25372 34552 25378 34604
rect 26237 34595 26295 34601
rect 26237 34561 26249 34595
rect 26283 34592 26295 34595
rect 26602 34592 26608 34604
rect 26283 34564 26608 34592
rect 26283 34561 26295 34564
rect 26237 34555 26295 34561
rect 26602 34552 26608 34564
rect 26660 34552 26666 34604
rect 26988 34601 27016 34632
rect 27338 34620 27344 34672
rect 27396 34660 27402 34672
rect 27396 34632 28764 34660
rect 27396 34620 27402 34632
rect 26973 34595 27031 34601
rect 26973 34561 26985 34595
rect 27019 34592 27031 34595
rect 27801 34595 27859 34601
rect 27801 34592 27813 34595
rect 27019 34564 27813 34592
rect 27019 34561 27031 34564
rect 26973 34555 27031 34561
rect 27801 34561 27813 34564
rect 27847 34561 27859 34595
rect 27801 34555 27859 34561
rect 28074 34552 28080 34604
rect 28132 34592 28138 34604
rect 28629 34595 28687 34601
rect 28629 34592 28641 34595
rect 28132 34564 28641 34592
rect 28132 34552 28138 34564
rect 28629 34561 28641 34564
rect 28675 34561 28687 34595
rect 28736 34592 28764 34632
rect 28994 34620 29000 34672
rect 29052 34660 29058 34672
rect 31205 34663 31263 34669
rect 29052 34632 29592 34660
rect 29052 34620 29058 34632
rect 29319 34595 29377 34601
rect 29319 34592 29331 34595
rect 28736 34564 29331 34592
rect 28629 34555 28687 34561
rect 29319 34561 29331 34564
rect 29365 34561 29377 34595
rect 29454 34592 29460 34604
rect 29415 34564 29460 34592
rect 29319 34555 29377 34561
rect 29454 34552 29460 34564
rect 29512 34552 29518 34604
rect 29564 34601 29592 34632
rect 31205 34629 31217 34663
rect 31251 34660 31263 34663
rect 32324 34660 32352 34688
rect 31251 34632 32352 34660
rect 36173 34663 36231 34669
rect 31251 34629 31263 34632
rect 31205 34623 31263 34629
rect 36173 34629 36185 34663
rect 36219 34660 36231 34663
rect 43438 34660 43444 34672
rect 36219 34632 43444 34660
rect 36219 34629 36231 34632
rect 36173 34623 36231 34629
rect 43438 34620 43444 34632
rect 43496 34620 43502 34672
rect 29549 34595 29607 34601
rect 29549 34561 29561 34595
rect 29595 34561 29607 34595
rect 29730 34592 29736 34604
rect 29691 34564 29736 34592
rect 29549 34555 29607 34561
rect 29730 34552 29736 34564
rect 29788 34552 29794 34604
rect 30098 34552 30104 34604
rect 30156 34592 30162 34604
rect 31389 34595 31447 34601
rect 31389 34592 31401 34595
rect 30156 34564 31401 34592
rect 30156 34552 30162 34564
rect 31389 34561 31401 34564
rect 31435 34561 31447 34595
rect 31389 34555 31447 34561
rect 31754 34552 31760 34604
rect 31812 34592 31818 34604
rect 32381 34595 32439 34601
rect 32381 34592 32393 34595
rect 31812 34564 32393 34592
rect 31812 34552 31818 34564
rect 32381 34561 32393 34564
rect 32427 34561 32439 34595
rect 32381 34555 32439 34561
rect 47302 34552 47308 34604
rect 47360 34592 47366 34604
rect 47581 34595 47639 34601
rect 47581 34592 47593 34595
rect 47360 34564 47593 34592
rect 47360 34552 47366 34564
rect 47581 34561 47593 34564
rect 47627 34561 47639 34595
rect 47581 34555 47639 34561
rect 23658 34524 23664 34536
rect 21744 34496 21864 34524
rect 15194 34416 15200 34468
rect 15252 34456 15258 34468
rect 16390 34456 16396 34468
rect 15252 34428 16396 34456
rect 15252 34416 15258 34428
rect 16390 34416 16396 34428
rect 16448 34416 16454 34468
rect 1394 34348 1400 34400
rect 1452 34388 1458 34400
rect 2041 34391 2099 34397
rect 2041 34388 2053 34391
rect 1452 34360 2053 34388
rect 1452 34348 1458 34360
rect 2041 34357 2053 34360
rect 2087 34357 2099 34391
rect 21836 34388 21864 34496
rect 22848 34496 23664 34524
rect 22848 34388 22876 34496
rect 23658 34484 23664 34496
rect 23716 34484 23722 34536
rect 23750 34484 23756 34536
rect 23808 34524 23814 34536
rect 23937 34527 23995 34533
rect 23937 34524 23949 34527
rect 23808 34496 23949 34524
rect 23808 34484 23814 34496
rect 23937 34493 23949 34496
rect 23983 34493 23995 34527
rect 23937 34487 23995 34493
rect 25593 34527 25651 34533
rect 25593 34493 25605 34527
rect 25639 34524 25651 34527
rect 26142 34524 26148 34536
rect 25639 34496 26148 34524
rect 25639 34493 25651 34496
rect 25593 34487 25651 34493
rect 26142 34484 26148 34496
rect 26200 34484 26206 34536
rect 29089 34527 29147 34533
rect 29089 34493 29101 34527
rect 29135 34524 29147 34527
rect 30374 34524 30380 34536
rect 29135 34496 30380 34524
rect 29135 34493 29147 34496
rect 29089 34487 29147 34493
rect 30374 34484 30380 34496
rect 30432 34484 30438 34536
rect 31573 34527 31631 34533
rect 31573 34493 31585 34527
rect 31619 34524 31631 34527
rect 31938 34524 31944 34536
rect 31619 34496 31944 34524
rect 31619 34493 31631 34496
rect 31573 34487 31631 34493
rect 31938 34484 31944 34496
rect 31996 34484 32002 34536
rect 32122 34524 32128 34536
rect 32083 34496 32128 34524
rect 32122 34484 32128 34496
rect 32180 34484 32186 34536
rect 33870 34484 33876 34536
rect 33928 34524 33934 34536
rect 34333 34527 34391 34533
rect 34333 34524 34345 34527
rect 33928 34496 34345 34524
rect 33928 34484 33934 34496
rect 34333 34493 34345 34496
rect 34379 34493 34391 34527
rect 34514 34524 34520 34536
rect 34475 34496 34520 34524
rect 34333 34487 34391 34493
rect 34514 34484 34520 34496
rect 34572 34484 34578 34536
rect 27157 34459 27215 34465
rect 27157 34425 27169 34459
rect 27203 34456 27215 34459
rect 27798 34456 27804 34468
rect 27203 34428 27804 34456
rect 27203 34425 27215 34428
rect 27157 34419 27215 34425
rect 27798 34416 27804 34428
rect 27856 34456 27862 34468
rect 28166 34456 28172 34468
rect 27856 34428 28172 34456
rect 27856 34416 27862 34428
rect 28166 34416 28172 34428
rect 28224 34416 28230 34468
rect 47026 34456 47032 34468
rect 46987 34428 47032 34456
rect 47026 34416 47032 34428
rect 47084 34416 47090 34468
rect 21836 34360 22876 34388
rect 2041 34351 2099 34357
rect 23474 34348 23480 34400
rect 23532 34388 23538 34400
rect 24949 34391 25007 34397
rect 24949 34388 24961 34391
rect 23532 34360 24961 34388
rect 23532 34348 23538 34360
rect 24949 34357 24961 34360
rect 24995 34357 25007 34391
rect 24949 34351 25007 34357
rect 25130 34348 25136 34400
rect 25188 34388 25194 34400
rect 25866 34388 25872 34400
rect 25188 34360 25872 34388
rect 25188 34348 25194 34360
rect 25866 34348 25872 34360
rect 25924 34348 25930 34400
rect 27893 34391 27951 34397
rect 27893 34357 27905 34391
rect 27939 34388 27951 34391
rect 28074 34388 28080 34400
rect 27939 34360 28080 34388
rect 27939 34357 27951 34360
rect 27893 34351 27951 34357
rect 28074 34348 28080 34360
rect 28132 34348 28138 34400
rect 28350 34348 28356 34400
rect 28408 34388 28414 34400
rect 28445 34391 28503 34397
rect 28445 34388 28457 34391
rect 28408 34360 28457 34388
rect 28408 34348 28414 34360
rect 28445 34357 28457 34360
rect 28491 34357 28503 34391
rect 28445 34351 28503 34357
rect 29178 34348 29184 34400
rect 29236 34388 29242 34400
rect 33502 34388 33508 34400
rect 29236 34360 33508 34388
rect 29236 34348 29242 34360
rect 33502 34348 33508 34360
rect 33560 34348 33566 34400
rect 46290 34348 46296 34400
rect 46348 34388 46354 34400
rect 46385 34391 46443 34397
rect 46385 34388 46397 34391
rect 46348 34360 46397 34388
rect 46348 34348 46354 34360
rect 46385 34357 46397 34360
rect 46431 34357 46443 34391
rect 47670 34388 47676 34400
rect 47631 34360 47676 34388
rect 46385 34351 46443 34357
rect 47670 34348 47676 34360
rect 47728 34348 47734 34400
rect 1104 34298 48852 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 48852 34298
rect 1104 34224 48852 34246
rect 13078 34144 13084 34196
rect 13136 34184 13142 34196
rect 16301 34187 16359 34193
rect 16301 34184 16313 34187
rect 13136 34156 16313 34184
rect 13136 34144 13142 34156
rect 16301 34153 16313 34156
rect 16347 34153 16359 34187
rect 16301 34147 16359 34153
rect 1394 34048 1400 34060
rect 1355 34020 1400 34048
rect 1394 34008 1400 34020
rect 1452 34008 1458 34060
rect 2774 34008 2780 34060
rect 2832 34048 2838 34060
rect 2832 34020 2877 34048
rect 2832 34008 2838 34020
rect 14921 33983 14979 33989
rect 14921 33949 14933 33983
rect 14967 33980 14979 33983
rect 15562 33980 15568 33992
rect 14967 33952 15568 33980
rect 14967 33949 14979 33952
rect 14921 33943 14979 33949
rect 15562 33940 15568 33952
rect 15620 33940 15626 33992
rect 16316 33980 16344 34147
rect 18138 34144 18144 34196
rect 18196 34184 18202 34196
rect 18693 34187 18751 34193
rect 18693 34184 18705 34187
rect 18196 34156 18705 34184
rect 18196 34144 18202 34156
rect 18693 34153 18705 34156
rect 18739 34153 18751 34187
rect 18693 34147 18751 34153
rect 22738 34144 22744 34196
rect 22796 34184 22802 34196
rect 24765 34187 24823 34193
rect 24765 34184 24777 34187
rect 22796 34156 24777 34184
rect 22796 34144 22802 34156
rect 24765 34153 24777 34156
rect 24811 34153 24823 34187
rect 24765 34147 24823 34153
rect 25225 34187 25283 34193
rect 25225 34153 25237 34187
rect 25271 34184 25283 34187
rect 25498 34184 25504 34196
rect 25271 34156 25504 34184
rect 25271 34153 25283 34156
rect 25225 34147 25283 34153
rect 25498 34144 25504 34156
rect 25556 34144 25562 34196
rect 25958 34184 25964 34196
rect 25919 34156 25964 34184
rect 25958 34144 25964 34156
rect 26016 34144 26022 34196
rect 26234 34184 26240 34196
rect 26195 34156 26240 34184
rect 26234 34144 26240 34156
rect 26292 34144 26298 34196
rect 28074 34144 28080 34196
rect 28132 34184 28138 34196
rect 31202 34184 31208 34196
rect 28132 34156 31208 34184
rect 28132 34144 28138 34156
rect 31202 34144 31208 34156
rect 31260 34144 31266 34196
rect 31389 34187 31447 34193
rect 31389 34153 31401 34187
rect 31435 34184 31447 34187
rect 31754 34184 31760 34196
rect 31435 34156 31760 34184
rect 31435 34153 31447 34156
rect 31389 34147 31447 34153
rect 31754 34144 31760 34156
rect 31812 34144 31818 34196
rect 34514 34144 34520 34196
rect 34572 34184 34578 34196
rect 34793 34187 34851 34193
rect 34793 34184 34805 34187
rect 34572 34156 34805 34184
rect 34572 34144 34578 34156
rect 34793 34153 34805 34156
rect 34839 34153 34851 34187
rect 34793 34147 34851 34153
rect 16390 34076 16396 34128
rect 16448 34116 16454 34128
rect 23934 34116 23940 34128
rect 16448 34088 23940 34116
rect 16448 34076 16454 34088
rect 23934 34076 23940 34088
rect 23992 34076 23998 34128
rect 26970 34116 26976 34128
rect 26931 34088 26976 34116
rect 26970 34076 26976 34088
rect 27028 34076 27034 34128
rect 47210 34116 47216 34128
rect 46308 34088 47216 34116
rect 21266 34008 21272 34060
rect 21324 34048 21330 34060
rect 24854 34048 24860 34060
rect 21324 34020 22094 34048
rect 24815 34020 24860 34048
rect 21324 34008 21330 34020
rect 16853 33983 16911 33989
rect 16853 33980 16865 33983
rect 16316 33952 16865 33980
rect 16853 33949 16865 33952
rect 16899 33949 16911 33983
rect 16853 33943 16911 33949
rect 18325 33983 18383 33989
rect 18325 33949 18337 33983
rect 18371 33980 18383 33983
rect 19242 33980 19248 33992
rect 18371 33952 19248 33980
rect 18371 33949 18383 33952
rect 18325 33943 18383 33949
rect 19242 33940 19248 33952
rect 19300 33940 19306 33992
rect 21361 33983 21419 33989
rect 21361 33949 21373 33983
rect 21407 33949 21419 33983
rect 21361 33943 21419 33949
rect 21637 33983 21695 33989
rect 21637 33949 21649 33983
rect 21683 33980 21695 33983
rect 21818 33980 21824 33992
rect 21683 33952 21824 33980
rect 21683 33949 21695 33952
rect 21637 33943 21695 33949
rect 1581 33915 1639 33921
rect 1581 33881 1593 33915
rect 1627 33912 1639 33915
rect 2130 33912 2136 33924
rect 1627 33884 2136 33912
rect 1627 33881 1639 33884
rect 1581 33875 1639 33881
rect 2130 33872 2136 33884
rect 2188 33872 2194 33924
rect 15188 33915 15246 33921
rect 15188 33881 15200 33915
rect 15234 33912 15246 33915
rect 15470 33912 15476 33924
rect 15234 33884 15476 33912
rect 15234 33881 15246 33884
rect 15188 33875 15246 33881
rect 15470 33872 15476 33884
rect 15528 33872 15534 33924
rect 16669 33915 16727 33921
rect 16669 33881 16681 33915
rect 16715 33912 16727 33915
rect 17494 33912 17500 33924
rect 16715 33884 17500 33912
rect 16715 33881 16727 33884
rect 16669 33875 16727 33881
rect 17494 33872 17500 33884
rect 17552 33872 17558 33924
rect 18509 33915 18567 33921
rect 18509 33881 18521 33915
rect 18555 33912 18567 33915
rect 19426 33912 19432 33924
rect 18555 33884 19432 33912
rect 18555 33881 18567 33884
rect 18509 33875 18567 33881
rect 19426 33872 19432 33884
rect 19484 33872 19490 33924
rect 21376 33912 21404 33943
rect 21818 33940 21824 33952
rect 21876 33940 21882 33992
rect 22066 33980 22094 34020
rect 24854 34008 24860 34020
rect 24912 34008 24918 34060
rect 26326 34048 26332 34060
rect 25884 34020 26332 34048
rect 25041 33983 25099 33989
rect 22066 33952 24900 33980
rect 22278 33912 22284 33924
rect 21376 33884 22284 33912
rect 22278 33872 22284 33884
rect 22336 33872 22342 33924
rect 23474 33912 23480 33924
rect 23435 33884 23480 33912
rect 23474 33872 23480 33884
rect 23532 33872 23538 33924
rect 23661 33915 23719 33921
rect 23661 33881 23673 33915
rect 23707 33912 23719 33915
rect 23750 33912 23756 33924
rect 23707 33884 23756 33912
rect 23707 33881 23719 33884
rect 23661 33875 23719 33881
rect 23750 33872 23756 33884
rect 23808 33872 23814 33924
rect 24670 33872 24676 33924
rect 24728 33912 24734 33924
rect 24765 33915 24823 33921
rect 24765 33912 24777 33915
rect 24728 33884 24777 33912
rect 24728 33872 24734 33884
rect 24765 33881 24777 33884
rect 24811 33881 24823 33915
rect 24872 33912 24900 33952
rect 25041 33949 25053 33983
rect 25087 33980 25099 33983
rect 25130 33980 25136 33992
rect 25087 33952 25136 33980
rect 25087 33949 25099 33952
rect 25041 33943 25099 33949
rect 25130 33940 25136 33952
rect 25188 33940 25194 33992
rect 25884 33989 25912 34020
rect 26326 34008 26332 34020
rect 26384 34008 26390 34060
rect 26602 34048 26608 34060
rect 26515 34020 26608 34048
rect 26602 34008 26608 34020
rect 26660 34048 26666 34060
rect 27525 34051 27583 34057
rect 27525 34048 27537 34051
rect 26660 34020 27537 34048
rect 26660 34008 26666 34020
rect 27525 34017 27537 34020
rect 27571 34017 27583 34051
rect 32398 34048 32404 34060
rect 27525 34011 27583 34017
rect 30944 34020 31800 34048
rect 25869 33983 25927 33989
rect 25869 33949 25881 33983
rect 25915 33949 25927 33983
rect 25869 33943 25927 33949
rect 26053 33983 26111 33989
rect 26053 33949 26065 33983
rect 26099 33980 26111 33983
rect 26620 33980 26648 34008
rect 26099 33952 26648 33980
rect 27433 33983 27491 33989
rect 26099 33949 26111 33952
rect 26053 33943 26111 33949
rect 27433 33949 27445 33983
rect 27479 33980 27491 33983
rect 27982 33980 27988 33992
rect 27479 33952 27988 33980
rect 27479 33949 27491 33952
rect 27433 33943 27491 33949
rect 26789 33915 26847 33921
rect 26789 33912 26801 33915
rect 24872 33884 26801 33912
rect 24765 33875 24823 33881
rect 26789 33881 26801 33884
rect 26835 33881 26847 33915
rect 26789 33875 26847 33881
rect 17034 33844 17040 33856
rect 16995 33816 17040 33844
rect 17034 33804 17040 33816
rect 17092 33804 17098 33856
rect 17126 33804 17132 33856
rect 17184 33844 17190 33856
rect 23566 33844 23572 33856
rect 17184 33816 23572 33844
rect 17184 33804 17190 33816
rect 23566 33804 23572 33816
rect 23624 33804 23630 33856
rect 23842 33844 23848 33856
rect 23803 33816 23848 33844
rect 23842 33804 23848 33816
rect 23900 33804 23906 33856
rect 24394 33804 24400 33856
rect 24452 33844 24458 33856
rect 27448 33844 27476 33943
rect 27982 33940 27988 33952
rect 28040 33940 28046 33992
rect 28350 33940 28356 33992
rect 28408 33980 28414 33992
rect 28813 33983 28871 33989
rect 28813 33980 28825 33983
rect 28408 33952 28825 33980
rect 28408 33940 28414 33952
rect 28813 33949 28825 33952
rect 28859 33949 28871 33983
rect 29546 33980 29552 33992
rect 29507 33952 29552 33980
rect 28813 33943 28871 33949
rect 29546 33940 29552 33952
rect 29604 33940 29610 33992
rect 28626 33912 28632 33924
rect 28587 33884 28632 33912
rect 28626 33872 28632 33884
rect 28684 33872 28690 33924
rect 29086 33872 29092 33924
rect 29144 33912 29150 33924
rect 29794 33915 29852 33921
rect 29794 33912 29806 33915
rect 29144 33884 29806 33912
rect 29144 33872 29150 33884
rect 29794 33881 29806 33884
rect 29840 33881 29852 33915
rect 29794 33875 29852 33881
rect 30944 33856 30972 34020
rect 31202 33940 31208 33992
rect 31260 33980 31266 33992
rect 31772 33989 31800 34020
rect 31864 34020 32404 34048
rect 31864 33989 31892 34020
rect 32398 34008 32404 34020
rect 32456 34008 32462 34060
rect 46308 34057 46336 34088
rect 47210 34076 47216 34088
rect 47268 34076 47274 34128
rect 46293 34051 46351 34057
rect 46293 34017 46305 34051
rect 46339 34017 46351 34051
rect 46293 34011 46351 34017
rect 46477 34051 46535 34057
rect 46477 34017 46489 34051
rect 46523 34048 46535 34051
rect 47670 34048 47676 34060
rect 46523 34020 47676 34048
rect 46523 34017 46535 34020
rect 46477 34011 46535 34017
rect 47670 34008 47676 34020
rect 47728 34008 47734 34060
rect 48130 34048 48136 34060
rect 48091 34020 48136 34048
rect 48130 34008 48136 34020
rect 48188 34008 48194 34060
rect 31665 33983 31723 33989
rect 31665 33980 31677 33983
rect 31260 33952 31677 33980
rect 31260 33940 31266 33952
rect 31665 33949 31677 33952
rect 31711 33949 31723 33983
rect 31665 33943 31723 33949
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33949 31815 33983
rect 31757 33943 31815 33949
rect 31849 33983 31907 33989
rect 31849 33949 31861 33983
rect 31895 33949 31907 33983
rect 31849 33943 31907 33949
rect 31938 33940 31944 33992
rect 31996 33980 32002 33992
rect 32033 33983 32091 33989
rect 32033 33980 32045 33983
rect 31996 33952 32045 33980
rect 31996 33940 32002 33952
rect 32033 33949 32045 33952
rect 32079 33949 32091 33983
rect 32033 33943 32091 33949
rect 32493 33983 32551 33989
rect 32493 33949 32505 33983
rect 32539 33949 32551 33983
rect 32493 33943 32551 33949
rect 32122 33912 32128 33924
rect 31772 33884 32128 33912
rect 31772 33856 31800 33884
rect 32122 33872 32128 33884
rect 32180 33912 32186 33924
rect 32508 33912 32536 33943
rect 33318 33940 33324 33992
rect 33376 33980 33382 33992
rect 33962 33980 33968 33992
rect 33376 33952 33968 33980
rect 33376 33940 33382 33952
rect 33962 33940 33968 33952
rect 34020 33980 34026 33992
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34020 33952 34713 33980
rect 34020 33940 34026 33952
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 32180 33884 32536 33912
rect 32180 33872 32186 33884
rect 32582 33872 32588 33924
rect 32640 33912 32646 33924
rect 32738 33915 32796 33921
rect 32738 33912 32750 33915
rect 32640 33884 32750 33912
rect 32640 33872 32646 33884
rect 32738 33881 32750 33884
rect 32784 33881 32796 33915
rect 32738 33875 32796 33881
rect 28994 33844 29000 33856
rect 24452 33816 27476 33844
rect 28955 33816 29000 33844
rect 24452 33804 24458 33816
rect 28994 33804 29000 33816
rect 29052 33804 29058 33856
rect 30926 33844 30932 33856
rect 30887 33816 30932 33844
rect 30926 33804 30932 33816
rect 30984 33804 30990 33856
rect 31754 33804 31760 33856
rect 31812 33804 31818 33856
rect 33870 33844 33876 33856
rect 33831 33816 33876 33844
rect 33870 33804 33876 33816
rect 33928 33804 33934 33856
rect 47946 33804 47952 33856
rect 48004 33844 48010 33856
rect 48130 33844 48136 33856
rect 48004 33816 48136 33844
rect 48004 33804 48010 33816
rect 48130 33804 48136 33816
rect 48188 33804 48194 33856
rect 1104 33754 48852 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 48852 33754
rect 1104 33680 48852 33702
rect 2130 33640 2136 33652
rect 2091 33612 2136 33640
rect 2130 33600 2136 33612
rect 2188 33600 2194 33652
rect 15470 33640 15476 33652
rect 15431 33612 15476 33640
rect 15470 33600 15476 33612
rect 15528 33600 15534 33652
rect 17954 33600 17960 33652
rect 18012 33640 18018 33652
rect 18509 33643 18567 33649
rect 18509 33640 18521 33643
rect 18012 33612 18521 33640
rect 18012 33600 18018 33612
rect 18509 33609 18521 33612
rect 18555 33609 18567 33643
rect 22370 33640 22376 33652
rect 22331 33612 22376 33640
rect 18509 33603 18567 33609
rect 22370 33600 22376 33612
rect 22428 33600 22434 33652
rect 23566 33600 23572 33652
rect 23624 33640 23630 33652
rect 24118 33640 24124 33652
rect 23624 33612 24124 33640
rect 23624 33600 23630 33612
rect 24118 33600 24124 33612
rect 24176 33600 24182 33652
rect 28626 33640 28632 33652
rect 28587 33612 28632 33640
rect 28626 33600 28632 33612
rect 28684 33600 28690 33652
rect 28997 33643 29055 33649
rect 28997 33609 29009 33643
rect 29043 33640 29055 33643
rect 30926 33640 30932 33652
rect 29043 33612 30932 33640
rect 29043 33609 29055 33612
rect 28997 33603 29055 33609
rect 30926 33600 30932 33612
rect 30984 33600 30990 33652
rect 32125 33643 32183 33649
rect 32125 33609 32137 33643
rect 32171 33640 32183 33643
rect 32582 33640 32588 33652
rect 32171 33612 32588 33640
rect 32171 33609 32183 33612
rect 32125 33603 32183 33609
rect 32582 33600 32588 33612
rect 32640 33600 32646 33652
rect 33410 33640 33416 33652
rect 33371 33612 33416 33640
rect 33410 33600 33416 33612
rect 33468 33600 33474 33652
rect 33502 33600 33508 33652
rect 33560 33640 33566 33652
rect 46017 33643 46075 33649
rect 33560 33612 45554 33640
rect 33560 33600 33566 33612
rect 17034 33572 17040 33584
rect 15948 33544 17040 33572
rect 2041 33507 2099 33513
rect 2041 33473 2053 33507
rect 2087 33504 2099 33507
rect 2222 33504 2228 33516
rect 2087 33476 2228 33504
rect 2087 33473 2099 33476
rect 2041 33467 2099 33473
rect 2222 33464 2228 33476
rect 2280 33464 2286 33516
rect 14366 33464 14372 33516
rect 14424 33504 14430 33516
rect 15948 33513 15976 33544
rect 17034 33532 17040 33544
rect 17092 33532 17098 33584
rect 17862 33572 17868 33584
rect 17328 33544 17868 33572
rect 15749 33507 15807 33513
rect 15749 33504 15761 33507
rect 14424 33476 15761 33504
rect 14424 33464 14430 33476
rect 15749 33473 15761 33476
rect 15795 33473 15807 33507
rect 15749 33467 15807 33473
rect 15841 33507 15899 33513
rect 15841 33473 15853 33507
rect 15887 33473 15899 33507
rect 15841 33467 15899 33473
rect 15933 33507 15991 33513
rect 15933 33473 15945 33507
rect 15979 33473 15991 33507
rect 15933 33467 15991 33473
rect 16117 33507 16175 33513
rect 16117 33473 16129 33507
rect 16163 33504 16175 33507
rect 17328 33504 17356 33544
rect 17862 33532 17868 33544
rect 17920 33532 17926 33584
rect 18417 33575 18475 33581
rect 18417 33541 18429 33575
rect 18463 33572 18475 33575
rect 21266 33572 21272 33584
rect 18463 33544 21272 33572
rect 18463 33541 18475 33544
rect 18417 33535 18475 33541
rect 21266 33532 21272 33544
rect 21324 33532 21330 33584
rect 22278 33572 22284 33584
rect 22239 33544 22284 33572
rect 22278 33532 22284 33544
rect 22336 33532 22342 33584
rect 25130 33532 25136 33584
rect 25188 33572 25194 33584
rect 25188 33544 25544 33572
rect 25188 33532 25194 33544
rect 17494 33504 17500 33516
rect 16163 33476 17356 33504
rect 17455 33476 17500 33504
rect 16163 33473 16175 33476
rect 16117 33467 16175 33473
rect 15856 33436 15884 33467
rect 17494 33464 17500 33476
rect 17552 33464 17558 33516
rect 17678 33504 17684 33516
rect 17639 33476 17684 33504
rect 17678 33464 17684 33476
rect 17736 33464 17742 33516
rect 19334 33464 19340 33516
rect 19392 33504 19398 33516
rect 19613 33507 19671 33513
rect 19613 33504 19625 33507
rect 19392 33476 19625 33504
rect 19392 33464 19398 33476
rect 19613 33473 19625 33476
rect 19659 33473 19671 33507
rect 19613 33467 19671 33473
rect 23566 33464 23572 33516
rect 23624 33507 23630 33516
rect 23661 33507 23719 33513
rect 23624 33479 23673 33507
rect 23624 33464 23630 33479
rect 23661 33473 23673 33479
rect 23707 33473 23719 33507
rect 23661 33467 23719 33473
rect 23753 33507 23811 33513
rect 23753 33473 23765 33507
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 17126 33436 17132 33448
rect 15856 33408 17132 33436
rect 17126 33396 17132 33408
rect 17184 33396 17190 33448
rect 17221 33439 17279 33445
rect 17221 33405 17233 33439
rect 17267 33436 17279 33439
rect 17696 33436 17724 33464
rect 17267 33408 17724 33436
rect 17267 33405 17279 33408
rect 17221 33399 17279 33405
rect 22094 33396 22100 33448
rect 22152 33436 22158 33448
rect 22462 33436 22468 33448
rect 22152 33408 22468 33436
rect 22152 33396 22158 33408
rect 22462 33396 22468 33408
rect 22520 33436 22526 33448
rect 23768 33436 23796 33467
rect 23842 33464 23848 33516
rect 23900 33504 23906 33516
rect 23900 33476 23945 33504
rect 23900 33464 23906 33476
rect 24026 33464 24032 33516
rect 24084 33504 24090 33516
rect 25406 33504 25412 33516
rect 24084 33476 24129 33504
rect 25367 33476 25412 33504
rect 24084 33464 24090 33476
rect 25406 33464 25412 33476
rect 25464 33464 25470 33516
rect 25516 33513 25544 33544
rect 27154 33532 27160 33584
rect 27212 33572 27218 33584
rect 27212 33544 29500 33572
rect 27212 33532 27218 33544
rect 25501 33507 25559 33513
rect 25501 33473 25513 33507
rect 25547 33473 25559 33507
rect 25501 33467 25559 33473
rect 25593 33507 25651 33513
rect 25593 33473 25605 33507
rect 25639 33504 25651 33507
rect 25777 33507 25835 33513
rect 25639 33476 25728 33504
rect 25639 33473 25651 33476
rect 25593 33467 25651 33473
rect 22520 33408 23796 33436
rect 22520 33396 22526 33408
rect 24302 33396 24308 33448
rect 24360 33436 24366 33448
rect 25700 33436 25728 33476
rect 25777 33473 25789 33507
rect 25823 33473 25835 33507
rect 25777 33467 25835 33473
rect 27801 33507 27859 33513
rect 27801 33473 27813 33507
rect 27847 33473 27859 33507
rect 27801 33467 27859 33473
rect 27985 33507 28043 33513
rect 27985 33473 27997 33507
rect 28031 33473 28043 33507
rect 27985 33467 28043 33473
rect 28169 33507 28227 33513
rect 28169 33473 28181 33507
rect 28215 33504 28227 33507
rect 28902 33504 28908 33516
rect 28215 33476 28908 33504
rect 28215 33473 28227 33476
rect 28169 33467 28227 33473
rect 24360 33408 25728 33436
rect 24360 33396 24366 33408
rect 19797 33371 19855 33377
rect 19797 33337 19809 33371
rect 19843 33368 19855 33371
rect 20438 33368 20444 33380
rect 19843 33340 20444 33368
rect 19843 33337 19855 33340
rect 19797 33331 19855 33337
rect 20438 33328 20444 33340
rect 20496 33368 20502 33380
rect 23474 33368 23480 33380
rect 20496 33340 23480 33368
rect 20496 33328 20502 33340
rect 23474 33328 23480 33340
rect 23532 33328 23538 33380
rect 25038 33328 25044 33380
rect 25096 33368 25102 33380
rect 25792 33368 25820 33467
rect 25096 33340 25820 33368
rect 27816 33368 27844 33467
rect 28000 33436 28028 33467
rect 28902 33464 28908 33476
rect 28960 33464 28966 33516
rect 29362 33504 29368 33516
rect 29012 33476 29368 33504
rect 28350 33436 28356 33448
rect 28000 33408 28356 33436
rect 28350 33396 28356 33408
rect 28408 33396 28414 33448
rect 29012 33368 29040 33476
rect 29362 33464 29368 33476
rect 29420 33464 29426 33516
rect 29472 33504 29500 33544
rect 29546 33532 29552 33584
rect 29604 33572 29610 33584
rect 31754 33572 31760 33584
rect 29604 33544 31760 33572
rect 29604 33532 29610 33544
rect 30116 33513 30144 33544
rect 31754 33532 31760 33544
rect 31812 33532 31818 33584
rect 40862 33572 40868 33584
rect 31864 33544 40868 33572
rect 30374 33513 30380 33516
rect 30101 33507 30159 33513
rect 29472 33476 29960 33504
rect 29089 33439 29147 33445
rect 29089 33405 29101 33439
rect 29135 33405 29147 33439
rect 29089 33399 29147 33405
rect 29181 33439 29239 33445
rect 29181 33405 29193 33439
rect 29227 33436 29239 33439
rect 29822 33436 29828 33448
rect 29227 33408 29828 33436
rect 29227 33405 29239 33408
rect 29181 33399 29239 33405
rect 27816 33340 29040 33368
rect 25096 33328 25102 33340
rect 2866 33300 2872 33312
rect 2827 33272 2872 33300
rect 2866 33260 2872 33272
rect 2924 33260 2930 33312
rect 17218 33260 17224 33312
rect 17276 33300 17282 33312
rect 17865 33303 17923 33309
rect 17865 33300 17877 33303
rect 17276 33272 17877 33300
rect 17276 33260 17282 33272
rect 17865 33269 17877 33272
rect 17911 33269 17923 33303
rect 17865 33263 17923 33269
rect 23385 33303 23443 33309
rect 23385 33269 23397 33303
rect 23431 33300 23443 33303
rect 24026 33300 24032 33312
rect 23431 33272 24032 33300
rect 23431 33269 23443 33272
rect 23385 33263 23443 33269
rect 24026 33260 24032 33272
rect 24084 33260 24090 33312
rect 25133 33303 25191 33309
rect 25133 33269 25145 33303
rect 25179 33300 25191 33303
rect 25866 33300 25872 33312
rect 25179 33272 25872 33300
rect 25179 33269 25191 33272
rect 25133 33263 25191 33269
rect 25866 33260 25872 33272
rect 25924 33260 25930 33312
rect 25958 33260 25964 33312
rect 26016 33300 26022 33312
rect 27154 33300 27160 33312
rect 26016 33272 27160 33300
rect 26016 33260 26022 33272
rect 27154 33260 27160 33272
rect 27212 33300 27218 33312
rect 29104 33300 29132 33399
rect 29822 33396 29828 33408
rect 29880 33396 29886 33448
rect 27212 33272 29132 33300
rect 29932 33300 29960 33476
rect 30101 33473 30113 33507
rect 30147 33473 30159 33507
rect 30368 33504 30380 33513
rect 30335 33476 30380 33504
rect 30101 33467 30159 33473
rect 30368 33467 30380 33476
rect 30374 33464 30380 33467
rect 30432 33464 30438 33516
rect 31864 33436 31892 33544
rect 40862 33532 40868 33544
rect 40920 33532 40926 33584
rect 45526 33572 45554 33612
rect 46017 33609 46029 33643
rect 46063 33640 46075 33643
rect 46474 33640 46480 33652
rect 46063 33612 46480 33640
rect 46063 33609 46075 33612
rect 46017 33603 46075 33609
rect 46474 33600 46480 33612
rect 46532 33600 46538 33652
rect 48133 33575 48191 33581
rect 48133 33572 48145 33575
rect 45526 33544 48145 33572
rect 48133 33541 48145 33544
rect 48179 33541 48191 33575
rect 48133 33535 48191 33541
rect 32401 33507 32459 33513
rect 32401 33504 32413 33507
rect 31128 33408 31892 33436
rect 31956 33476 32413 33504
rect 31128 33300 31156 33408
rect 31202 33328 31208 33380
rect 31260 33368 31266 33380
rect 31956 33368 31984 33476
rect 32401 33473 32413 33476
rect 32447 33473 32459 33507
rect 32401 33467 32459 33473
rect 32493 33507 32551 33513
rect 32493 33473 32505 33507
rect 32539 33473 32551 33507
rect 32493 33467 32551 33473
rect 31260 33340 31984 33368
rect 31260 33328 31266 33340
rect 31478 33300 31484 33312
rect 29932 33272 31156 33300
rect 31439 33272 31484 33300
rect 27212 33260 27218 33272
rect 31478 33260 31484 33272
rect 31536 33300 31542 33312
rect 32508 33300 32536 33467
rect 32582 33464 32588 33516
rect 32640 33504 32646 33516
rect 32766 33504 32772 33516
rect 32640 33476 32685 33504
rect 32727 33476 32772 33504
rect 32640 33464 32646 33476
rect 32766 33464 32772 33476
rect 32824 33464 32830 33516
rect 33318 33504 33324 33516
rect 33279 33476 33324 33504
rect 33318 33464 33324 33476
rect 33376 33464 33382 33516
rect 45922 33504 45928 33516
rect 45883 33476 45928 33504
rect 45922 33464 45928 33476
rect 45980 33464 45986 33516
rect 46566 33504 46572 33516
rect 46527 33476 46572 33504
rect 46566 33464 46572 33476
rect 46624 33464 46630 33516
rect 47946 33504 47952 33516
rect 47907 33476 47952 33504
rect 47946 33464 47952 33476
rect 48004 33464 48010 33516
rect 31536 33272 32536 33300
rect 31536 33260 31542 33272
rect 46474 33260 46480 33312
rect 46532 33300 46538 33312
rect 46661 33303 46719 33309
rect 46661 33300 46673 33303
rect 46532 33272 46673 33300
rect 46532 33260 46538 33272
rect 46661 33269 46673 33272
rect 46707 33269 46719 33303
rect 46661 33263 46719 33269
rect 47946 33260 47952 33312
rect 48004 33300 48010 33312
rect 48314 33300 48320 33312
rect 48004 33272 48320 33300
rect 48004 33260 48010 33272
rect 48314 33260 48320 33272
rect 48372 33260 48378 33312
rect 1104 33210 48852 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 48852 33210
rect 1104 33136 48852 33158
rect 13449 33099 13507 33105
rect 13449 33065 13461 33099
rect 13495 33096 13507 33099
rect 23566 33096 23572 33108
rect 13495 33068 14596 33096
rect 13495 33065 13507 33068
rect 13449 33059 13507 33065
rect 13906 33028 13912 33040
rect 13648 33000 13912 33028
rect 13262 32960 13268 32972
rect 13223 32932 13268 32960
rect 13262 32920 13268 32932
rect 13320 32920 13326 32972
rect 1762 32852 1768 32904
rect 1820 32892 1826 32904
rect 2590 32892 2596 32904
rect 1820 32864 2596 32892
rect 1820 32852 1826 32864
rect 2590 32852 2596 32864
rect 2648 32852 2654 32904
rect 2961 32895 3019 32901
rect 2961 32861 2973 32895
rect 3007 32892 3019 32895
rect 3970 32892 3976 32904
rect 3007 32864 3976 32892
rect 3007 32861 3019 32864
rect 2961 32855 3019 32861
rect 3970 32852 3976 32864
rect 4028 32852 4034 32904
rect 13173 32895 13231 32901
rect 13173 32861 13185 32895
rect 13219 32892 13231 32895
rect 13648 32892 13676 33000
rect 13906 32988 13912 33000
rect 13964 32988 13970 33040
rect 13219 32864 13676 32892
rect 13219 32861 13231 32864
rect 13173 32855 13231 32861
rect 13814 32852 13820 32904
rect 13872 32892 13878 32904
rect 14568 32901 14596 33068
rect 23216 33068 23572 33096
rect 17678 32988 17684 33040
rect 17736 33028 17742 33040
rect 17773 33031 17831 33037
rect 17773 33028 17785 33031
rect 17736 33000 17785 33028
rect 17736 32988 17742 33000
rect 17773 32997 17785 33000
rect 17819 33028 17831 33031
rect 17819 33000 20944 33028
rect 17819 32997 17831 33000
rect 17773 32991 17831 32997
rect 15562 32920 15568 32972
rect 15620 32960 15626 32972
rect 16393 32963 16451 32969
rect 16393 32960 16405 32963
rect 15620 32932 16405 32960
rect 15620 32920 15626 32932
rect 16393 32929 16405 32932
rect 16439 32929 16451 32963
rect 20806 32960 20812 32972
rect 16393 32923 16451 32929
rect 20088 32932 20812 32960
rect 14323 32895 14381 32901
rect 14553 32895 14611 32901
rect 14323 32892 14335 32895
rect 13872 32864 14335 32892
rect 13872 32852 13878 32864
rect 14323 32861 14335 32864
rect 14369 32861 14381 32895
rect 14323 32855 14381 32861
rect 14458 32889 14516 32895
rect 14458 32855 14470 32889
rect 14504 32855 14516 32889
rect 14553 32861 14565 32895
rect 14599 32861 14611 32895
rect 14734 32892 14740 32904
rect 14695 32864 14740 32892
rect 14553 32855 14611 32861
rect 14458 32849 14516 32855
rect 14734 32852 14740 32864
rect 14792 32852 14798 32904
rect 16942 32852 16948 32904
rect 17000 32892 17006 32904
rect 18138 32892 18144 32904
rect 17000 32864 18144 32892
rect 17000 32852 17006 32864
rect 18138 32852 18144 32864
rect 18196 32892 18202 32904
rect 18509 32895 18567 32901
rect 18509 32892 18521 32895
rect 18196 32864 18521 32892
rect 18196 32852 18202 32864
rect 18509 32861 18521 32864
rect 18555 32861 18567 32895
rect 18509 32855 18567 32861
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 20088 32901 20116 32932
rect 20806 32920 20812 32932
rect 20864 32920 20870 32972
rect 19889 32895 19947 32901
rect 19889 32892 19901 32895
rect 19208 32864 19901 32892
rect 19208 32852 19214 32864
rect 19889 32861 19901 32864
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 19981 32895 20039 32901
rect 19981 32861 19993 32895
rect 20027 32861 20039 32895
rect 19981 32855 20039 32861
rect 20073 32895 20131 32901
rect 20073 32861 20085 32895
rect 20119 32861 20131 32895
rect 20073 32855 20131 32861
rect 20257 32895 20315 32901
rect 20257 32861 20269 32895
rect 20303 32892 20315 32895
rect 20438 32892 20444 32904
rect 20303 32864 20444 32892
rect 20303 32861 20315 32864
rect 20257 32855 20315 32861
rect 14476 32768 14504 32849
rect 16666 32833 16672 32836
rect 16660 32787 16672 32833
rect 16724 32824 16730 32836
rect 18693 32827 18751 32833
rect 16724 32796 16760 32824
rect 16666 32784 16672 32787
rect 16724 32784 16730 32796
rect 18693 32793 18705 32827
rect 18739 32824 18751 32827
rect 19426 32824 19432 32836
rect 18739 32796 19432 32824
rect 18739 32793 18751 32796
rect 18693 32787 18751 32793
rect 19426 32784 19432 32796
rect 19484 32784 19490 32836
rect 19996 32824 20024 32855
rect 20438 32852 20444 32864
rect 20496 32852 20502 32904
rect 20916 32892 20944 33000
rect 21361 32963 21419 32969
rect 21361 32929 21373 32963
rect 21407 32960 21419 32963
rect 21818 32960 21824 32972
rect 21407 32932 21824 32960
rect 21407 32929 21419 32932
rect 21361 32923 21419 32929
rect 21818 32920 21824 32932
rect 21876 32960 21882 32972
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 21876 32932 22937 32960
rect 21876 32920 21882 32932
rect 22925 32929 22937 32932
rect 22971 32960 22983 32963
rect 23216 32960 23244 33068
rect 23566 33056 23572 33068
rect 23624 33056 23630 33108
rect 23845 33099 23903 33105
rect 23845 33065 23857 33099
rect 23891 33096 23903 33099
rect 24302 33096 24308 33108
rect 23891 33068 24308 33096
rect 23891 33065 23903 33068
rect 23845 33059 23903 33065
rect 24302 33056 24308 33068
rect 24360 33056 24366 33108
rect 32585 33099 32643 33105
rect 24964 33068 31754 33096
rect 24964 33028 24992 33068
rect 27154 33028 27160 33040
rect 22971 32932 23244 32960
rect 23308 33000 24992 33028
rect 27115 33000 27160 33028
rect 22971 32929 22983 32932
rect 22925 32923 22983 32929
rect 23308 32892 23336 33000
rect 27154 32988 27160 33000
rect 27212 32988 27218 33040
rect 28353 33031 28411 33037
rect 28353 32997 28365 33031
rect 28399 33028 28411 33031
rect 29086 33028 29092 33040
rect 28399 33000 29092 33028
rect 28399 32997 28411 33000
rect 28353 32991 28411 32997
rect 29086 32988 29092 33000
rect 29144 32988 29150 33040
rect 29362 32988 29368 33040
rect 29420 33028 29426 33040
rect 29549 33031 29607 33037
rect 29549 33028 29561 33031
rect 29420 33000 29561 33028
rect 29420 32988 29426 33000
rect 29549 32997 29561 33000
rect 29595 32997 29607 33031
rect 31726 33028 31754 33068
rect 32585 33065 32597 33099
rect 32631 33096 32643 33099
rect 32766 33096 32772 33108
rect 32631 33068 32772 33096
rect 32631 33065 32643 33068
rect 32585 33059 32643 33065
rect 32766 33056 32772 33068
rect 32824 33056 32830 33108
rect 31726 33000 35204 33028
rect 29549 32991 29607 32997
rect 23566 32920 23572 32972
rect 23624 32960 23630 32972
rect 24302 32960 24308 32972
rect 23624 32932 24308 32960
rect 23624 32920 23630 32932
rect 24302 32920 24308 32932
rect 24360 32960 24366 32972
rect 24360 32932 24624 32960
rect 24360 32920 24366 32932
rect 20916 32864 23336 32892
rect 23477 32895 23535 32901
rect 23477 32861 23489 32895
rect 23523 32892 23535 32895
rect 24596 32892 24624 32932
rect 24670 32920 24676 32972
rect 24728 32960 24734 32972
rect 24857 32963 24915 32969
rect 24857 32960 24869 32963
rect 24728 32932 24869 32960
rect 24728 32920 24734 32932
rect 24857 32929 24869 32932
rect 24903 32929 24915 32963
rect 24857 32923 24915 32929
rect 24949 32963 25007 32969
rect 24949 32929 24961 32963
rect 24995 32929 25007 32963
rect 24949 32923 25007 32929
rect 24964 32892 24992 32923
rect 29822 32920 29828 32972
rect 29880 32960 29886 32972
rect 35176 32969 35204 33000
rect 30101 32963 30159 32969
rect 30101 32960 30113 32963
rect 29880 32932 30113 32960
rect 29880 32920 29886 32932
rect 30101 32929 30113 32932
rect 30147 32929 30159 32963
rect 30101 32923 30159 32929
rect 35161 32963 35219 32969
rect 35161 32929 35173 32963
rect 35207 32929 35219 32963
rect 36998 32960 37004 32972
rect 36959 32932 37004 32960
rect 35161 32923 35219 32929
rect 36998 32920 37004 32932
rect 37056 32920 37062 32972
rect 46290 32960 46296 32972
rect 46251 32932 46296 32960
rect 46290 32920 46296 32932
rect 46348 32920 46354 32972
rect 46474 32960 46480 32972
rect 46435 32932 46480 32960
rect 46474 32920 46480 32932
rect 46532 32920 46538 32972
rect 48038 32960 48044 32972
rect 47999 32932 48044 32960
rect 48038 32920 48044 32932
rect 48096 32920 48102 32972
rect 25774 32892 25780 32904
rect 23523 32864 24440 32892
rect 24596 32864 24992 32892
rect 25735 32864 25780 32892
rect 23523 32861 23535 32864
rect 23477 32855 23535 32861
rect 20162 32824 20168 32836
rect 19996 32796 20168 32824
rect 20162 32784 20168 32796
rect 20220 32784 20226 32836
rect 21177 32827 21235 32833
rect 21177 32793 21189 32827
rect 21223 32824 21235 32827
rect 22002 32824 22008 32836
rect 21223 32796 22008 32824
rect 21223 32793 21235 32796
rect 21177 32787 21235 32793
rect 22002 32784 22008 32796
rect 22060 32784 22066 32836
rect 22649 32827 22707 32833
rect 22649 32793 22661 32827
rect 22695 32824 22707 32827
rect 22922 32824 22928 32836
rect 22695 32796 22928 32824
rect 22695 32793 22707 32796
rect 22649 32787 22707 32793
rect 22922 32784 22928 32796
rect 22980 32784 22986 32836
rect 23290 32784 23296 32836
rect 23348 32824 23354 32836
rect 23661 32827 23719 32833
rect 23661 32824 23673 32827
rect 23348 32796 23673 32824
rect 23348 32784 23354 32796
rect 23661 32793 23673 32796
rect 23707 32793 23719 32827
rect 23661 32787 23719 32793
rect 1762 32716 1768 32768
rect 1820 32756 1826 32768
rect 1857 32759 1915 32765
rect 1857 32756 1869 32759
rect 1820 32728 1869 32756
rect 1820 32716 1826 32728
rect 1857 32725 1869 32728
rect 1903 32725 1915 32759
rect 3050 32756 3056 32768
rect 3011 32728 3056 32756
rect 1857 32719 1915 32725
rect 3050 32716 3056 32728
rect 3108 32716 3114 32768
rect 14090 32756 14096 32768
rect 14051 32728 14096 32756
rect 14090 32716 14096 32728
rect 14148 32716 14154 32768
rect 14458 32716 14464 32768
rect 14516 32716 14522 32768
rect 19613 32759 19671 32765
rect 19613 32725 19625 32759
rect 19659 32756 19671 32759
rect 19978 32756 19984 32768
rect 19659 32728 19984 32756
rect 19659 32725 19671 32728
rect 19613 32719 19671 32725
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20714 32756 20720 32768
rect 20675 32728 20720 32756
rect 20714 32716 20720 32728
rect 20772 32716 20778 32768
rect 21082 32756 21088 32768
rect 21043 32728 21088 32756
rect 21082 32716 21088 32728
rect 21140 32716 21146 32768
rect 22186 32716 22192 32768
rect 22244 32756 22250 32768
rect 22281 32759 22339 32765
rect 22281 32756 22293 32759
rect 22244 32728 22293 32756
rect 22244 32716 22250 32728
rect 22281 32725 22293 32728
rect 22327 32725 22339 32759
rect 22281 32719 22339 32725
rect 22741 32759 22799 32765
rect 22741 32725 22753 32759
rect 22787 32756 22799 32759
rect 23106 32756 23112 32768
rect 22787 32728 23112 32756
rect 22787 32725 22799 32728
rect 22741 32719 22799 32725
rect 23106 32716 23112 32728
rect 23164 32716 23170 32768
rect 24412 32765 24440 32864
rect 25774 32852 25780 32864
rect 25832 32852 25838 32904
rect 25866 32852 25872 32904
rect 25924 32892 25930 32904
rect 26033 32895 26091 32901
rect 26033 32892 26045 32895
rect 25924 32864 26045 32892
rect 25924 32852 25930 32864
rect 26033 32861 26045 32864
rect 26079 32861 26091 32895
rect 26033 32855 26091 32861
rect 26970 32852 26976 32904
rect 27028 32892 27034 32904
rect 27709 32895 27767 32901
rect 27709 32892 27721 32895
rect 27028 32864 27721 32892
rect 27028 32852 27034 32864
rect 27709 32861 27721 32864
rect 27755 32861 27767 32895
rect 27709 32855 27767 32861
rect 28534 32852 28540 32904
rect 28592 32892 28598 32904
rect 28629 32895 28687 32901
rect 28629 32892 28641 32895
rect 28592 32864 28641 32892
rect 28592 32852 28598 32864
rect 28629 32861 28641 32864
rect 28675 32861 28687 32895
rect 28629 32855 28687 32861
rect 28721 32895 28779 32901
rect 28721 32861 28733 32895
rect 28767 32861 28779 32895
rect 28721 32855 28779 32861
rect 28813 32895 28871 32901
rect 28813 32861 28825 32895
rect 28859 32892 28871 32895
rect 28902 32892 28908 32904
rect 28859 32864 28908 32892
rect 28859 32861 28871 32864
rect 28813 32855 28871 32861
rect 27890 32824 27896 32836
rect 27851 32796 27896 32824
rect 27890 32784 27896 32796
rect 27948 32784 27954 32836
rect 28736 32824 28764 32855
rect 28902 32852 28908 32864
rect 28960 32852 28966 32904
rect 28994 32852 29000 32904
rect 29052 32892 29058 32904
rect 29730 32892 29736 32904
rect 29052 32864 29736 32892
rect 29052 32852 29058 32864
rect 29730 32852 29736 32864
rect 29788 32852 29794 32904
rect 29917 32895 29975 32901
rect 29917 32861 29929 32895
rect 29963 32892 29975 32895
rect 31478 32892 31484 32904
rect 29963 32864 31484 32892
rect 29963 32861 29975 32864
rect 29917 32855 29975 32861
rect 31478 32852 31484 32864
rect 31536 32852 31542 32904
rect 32217 32895 32275 32901
rect 32217 32861 32229 32895
rect 32263 32892 32275 32895
rect 33870 32892 33876 32904
rect 32263 32864 33876 32892
rect 32263 32861 32275 32864
rect 32217 32855 32275 32861
rect 33870 32852 33876 32864
rect 33928 32852 33934 32904
rect 29178 32824 29184 32836
rect 28736 32796 29184 32824
rect 29178 32784 29184 32796
rect 29236 32824 29242 32836
rect 29454 32824 29460 32836
rect 29236 32796 29460 32824
rect 29236 32784 29242 32796
rect 29454 32784 29460 32796
rect 29512 32784 29518 32836
rect 29748 32824 29776 32852
rect 30282 32824 30288 32836
rect 29748 32796 30288 32824
rect 30282 32784 30288 32796
rect 30340 32784 30346 32836
rect 32398 32824 32404 32836
rect 32359 32796 32404 32824
rect 32398 32784 32404 32796
rect 32456 32784 32462 32836
rect 35342 32824 35348 32836
rect 35303 32796 35348 32824
rect 35342 32784 35348 32796
rect 35400 32784 35406 32836
rect 24397 32759 24455 32765
rect 24397 32725 24409 32759
rect 24443 32725 24455 32759
rect 24397 32719 24455 32725
rect 24765 32759 24823 32765
rect 24765 32725 24777 32759
rect 24811 32756 24823 32759
rect 25958 32756 25964 32768
rect 24811 32728 25964 32756
rect 24811 32725 24823 32728
rect 24765 32719 24823 32725
rect 25958 32716 25964 32728
rect 26016 32716 26022 32768
rect 30006 32756 30012 32768
rect 29967 32728 30012 32756
rect 30006 32716 30012 32728
rect 30064 32716 30070 32768
rect 1104 32666 48852 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 48852 32666
rect 1104 32592 48852 32614
rect 10962 32512 10968 32564
rect 11020 32552 11026 32564
rect 12897 32555 12955 32561
rect 12897 32552 12909 32555
rect 11020 32524 12909 32552
rect 11020 32512 11026 32524
rect 12897 32521 12909 32524
rect 12943 32521 12955 32555
rect 12897 32515 12955 32521
rect 13262 32512 13268 32564
rect 13320 32552 13326 32564
rect 13633 32555 13691 32561
rect 13633 32552 13645 32555
rect 13320 32524 13645 32552
rect 13320 32512 13326 32524
rect 13633 32521 13645 32524
rect 13679 32521 13691 32555
rect 16666 32552 16672 32564
rect 16627 32524 16672 32552
rect 13633 32515 13691 32521
rect 16666 32512 16672 32524
rect 16724 32512 16730 32564
rect 17862 32512 17868 32564
rect 17920 32512 17926 32564
rect 20993 32555 21051 32561
rect 20993 32521 21005 32555
rect 21039 32552 21051 32555
rect 21082 32552 21088 32564
rect 21039 32524 21088 32552
rect 21039 32521 21051 32524
rect 20993 32515 21051 32521
rect 21082 32512 21088 32524
rect 21140 32552 21146 32564
rect 24946 32552 24952 32564
rect 21140 32524 24952 32552
rect 21140 32512 21146 32524
rect 24946 32512 24952 32524
rect 25004 32512 25010 32564
rect 25314 32552 25320 32564
rect 25275 32524 25320 32552
rect 25314 32512 25320 32524
rect 25372 32512 25378 32564
rect 26326 32552 26332 32564
rect 26287 32524 26332 32552
rect 26326 32512 26332 32524
rect 26384 32512 26390 32564
rect 30006 32552 30012 32564
rect 27816 32524 30012 32552
rect 14090 32444 14096 32496
rect 14148 32484 14154 32496
rect 14430 32487 14488 32493
rect 14430 32484 14442 32487
rect 14148 32456 14442 32484
rect 14148 32444 14154 32456
rect 14430 32453 14442 32456
rect 14476 32453 14488 32487
rect 17586 32484 17592 32496
rect 14430 32447 14488 32453
rect 17328 32456 17592 32484
rect 1762 32416 1768 32428
rect 1723 32388 1768 32416
rect 1762 32376 1768 32388
rect 1820 32376 1826 32428
rect 10870 32376 10876 32428
rect 10928 32416 10934 32428
rect 11773 32419 11831 32425
rect 11773 32416 11785 32419
rect 10928 32388 11785 32416
rect 10928 32376 10934 32388
rect 11773 32385 11785 32388
rect 11819 32385 11831 32419
rect 11773 32379 11831 32385
rect 13541 32419 13599 32425
rect 13541 32385 13553 32419
rect 13587 32385 13599 32419
rect 13541 32379 13599 32385
rect 13725 32419 13783 32425
rect 13725 32385 13737 32419
rect 13771 32416 13783 32419
rect 14274 32416 14280 32428
rect 13771 32388 14280 32416
rect 13771 32385 13783 32388
rect 13725 32379 13783 32385
rect 1946 32348 1952 32360
rect 1907 32320 1952 32348
rect 1946 32308 1952 32320
rect 2004 32308 2010 32360
rect 2774 32308 2780 32360
rect 2832 32348 2838 32360
rect 11517 32351 11575 32357
rect 2832 32320 2877 32348
rect 2832 32308 2838 32320
rect 11517 32317 11529 32351
rect 11563 32317 11575 32351
rect 13556 32348 13584 32379
rect 14274 32376 14280 32388
rect 14332 32376 14338 32428
rect 16574 32376 16580 32428
rect 16632 32416 16638 32428
rect 16945 32419 17003 32425
rect 16945 32416 16957 32419
rect 16632 32388 16957 32416
rect 16632 32376 16638 32388
rect 16945 32385 16957 32388
rect 16991 32385 17003 32419
rect 16945 32379 17003 32385
rect 17034 32419 17092 32425
rect 17034 32385 17046 32419
rect 17080 32385 17092 32419
rect 17034 32379 17092 32385
rect 17129 32422 17187 32428
rect 17129 32388 17141 32422
rect 17175 32416 17187 32422
rect 17218 32416 17224 32428
rect 17175 32388 17224 32416
rect 17129 32382 17187 32388
rect 13998 32348 14004 32360
rect 13556 32320 14004 32348
rect 11517 32311 11575 32317
rect 11532 32212 11560 32311
rect 13998 32308 14004 32320
rect 14056 32308 14062 32360
rect 14185 32351 14243 32357
rect 14185 32317 14197 32351
rect 14231 32317 14243 32351
rect 17049 32348 17077 32379
rect 17218 32376 17224 32388
rect 17276 32376 17282 32428
rect 17328 32425 17356 32456
rect 17586 32444 17592 32456
rect 17644 32484 17650 32496
rect 17880 32484 17908 32512
rect 18138 32484 18144 32496
rect 17644 32456 17908 32484
rect 18099 32456 18144 32484
rect 17644 32444 17650 32456
rect 18138 32444 18144 32456
rect 18196 32444 18202 32496
rect 20622 32484 20628 32496
rect 19628 32456 20628 32484
rect 17313 32419 17371 32425
rect 17313 32385 17325 32419
rect 17359 32385 17371 32419
rect 17862 32416 17868 32428
rect 17823 32388 17868 32416
rect 17313 32379 17371 32385
rect 17862 32376 17868 32388
rect 17920 32376 17926 32428
rect 18046 32416 18052 32428
rect 18007 32388 18052 32416
rect 18046 32376 18052 32388
rect 18104 32376 18110 32428
rect 19628 32425 19656 32456
rect 20622 32444 20628 32456
rect 20680 32484 20686 32496
rect 20680 32456 21864 32484
rect 20680 32444 20686 32456
rect 19886 32425 19892 32428
rect 19613 32419 19671 32425
rect 19613 32385 19625 32419
rect 19659 32385 19671 32419
rect 19880 32416 19892 32425
rect 19847 32388 19892 32416
rect 19613 32379 19671 32385
rect 19880 32379 19892 32388
rect 19886 32376 19892 32379
rect 19944 32376 19950 32428
rect 21836 32425 21864 32456
rect 22278 32444 22284 32496
rect 22336 32484 22342 32496
rect 23842 32484 23848 32496
rect 22336 32456 23848 32484
rect 22336 32444 22342 32456
rect 23842 32444 23848 32456
rect 23900 32444 23906 32496
rect 25774 32484 25780 32496
rect 23952 32456 24348 32484
rect 21821 32419 21879 32425
rect 21821 32385 21833 32419
rect 21867 32385 21879 32419
rect 21821 32379 21879 32385
rect 21910 32376 21916 32428
rect 21968 32416 21974 32428
rect 23952 32425 23980 32456
rect 22077 32419 22135 32425
rect 22077 32416 22089 32419
rect 21968 32388 22089 32416
rect 21968 32376 21974 32388
rect 22077 32385 22089 32388
rect 22123 32385 22135 32419
rect 22077 32379 22135 32385
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 23937 32379 23995 32385
rect 24026 32376 24032 32428
rect 24084 32416 24090 32428
rect 24193 32419 24251 32425
rect 24193 32416 24205 32419
rect 24084 32388 24205 32416
rect 24084 32376 24090 32388
rect 24193 32385 24205 32388
rect 24239 32385 24251 32419
rect 24320 32416 24348 32456
rect 25240 32456 25780 32484
rect 25240 32416 25268 32456
rect 25774 32444 25780 32456
rect 25832 32444 25838 32496
rect 24320 32388 25268 32416
rect 24193 32379 24251 32385
rect 25682 32376 25688 32428
rect 25740 32416 25746 32428
rect 25869 32419 25927 32425
rect 25869 32416 25881 32419
rect 25740 32388 25881 32416
rect 25740 32376 25746 32388
rect 25869 32385 25881 32388
rect 25915 32385 25927 32419
rect 26145 32419 26203 32425
rect 26145 32416 26157 32419
rect 25869 32379 25927 32385
rect 25976 32388 26157 32416
rect 17049 32320 17172 32348
rect 14185 32311 14243 32317
rect 14200 32280 14228 32311
rect 17144 32292 17172 32320
rect 24946 32308 24952 32360
rect 25004 32348 25010 32360
rect 25976 32348 26004 32388
rect 26145 32385 26157 32388
rect 26191 32385 26203 32419
rect 26145 32379 26203 32385
rect 25004 32320 26004 32348
rect 26053 32351 26111 32357
rect 25004 32308 25010 32320
rect 26053 32317 26065 32351
rect 26099 32317 26111 32351
rect 26160 32348 26188 32379
rect 26234 32376 26240 32428
rect 26292 32416 26298 32428
rect 27709 32419 27767 32425
rect 27709 32416 27721 32419
rect 26292 32388 27721 32416
rect 26292 32376 26298 32388
rect 27709 32385 27721 32388
rect 27755 32385 27767 32419
rect 27709 32379 27767 32385
rect 27338 32348 27344 32360
rect 26160 32320 27344 32348
rect 26053 32311 26111 32317
rect 12820 32252 14228 32280
rect 12710 32212 12716 32224
rect 11532 32184 12716 32212
rect 12710 32172 12716 32184
rect 12768 32212 12774 32224
rect 12820 32212 12848 32252
rect 17126 32240 17132 32292
rect 17184 32240 17190 32292
rect 26068 32280 26096 32311
rect 27338 32308 27344 32320
rect 27396 32308 27402 32360
rect 27816 32280 27844 32524
rect 30006 32512 30012 32524
rect 30064 32512 30070 32564
rect 27890 32444 27896 32496
rect 27948 32484 27954 32496
rect 30469 32487 30527 32493
rect 30469 32484 30481 32487
rect 27948 32456 30481 32484
rect 27948 32444 27954 32456
rect 30469 32453 30481 32456
rect 30515 32453 30527 32487
rect 30469 32447 30527 32453
rect 32217 32487 32275 32493
rect 32217 32453 32229 32487
rect 32263 32484 32275 32487
rect 33870 32484 33876 32496
rect 32263 32456 33876 32484
rect 32263 32453 32275 32456
rect 32217 32447 32275 32453
rect 33870 32444 33876 32456
rect 33928 32444 33934 32496
rect 28353 32419 28411 32425
rect 28353 32385 28365 32419
rect 28399 32385 28411 32419
rect 28353 32379 28411 32385
rect 28368 32348 28396 32379
rect 28442 32376 28448 32428
rect 28500 32416 28506 32428
rect 28537 32419 28595 32425
rect 28537 32416 28549 32419
rect 28500 32388 28549 32416
rect 28500 32376 28506 32388
rect 28537 32385 28549 32388
rect 28583 32385 28595 32419
rect 28537 32379 28595 32385
rect 28626 32376 28632 32428
rect 28684 32416 28690 32428
rect 28994 32416 29000 32428
rect 28684 32388 29000 32416
rect 28684 32376 28690 32388
rect 28994 32376 29000 32388
rect 29052 32376 29058 32428
rect 29549 32419 29607 32425
rect 29549 32385 29561 32419
rect 29595 32416 29607 32419
rect 31846 32416 31852 32428
rect 29595 32388 31852 32416
rect 29595 32385 29607 32388
rect 29549 32379 29607 32385
rect 31846 32376 31852 32388
rect 31904 32376 31910 32428
rect 32398 32416 32404 32428
rect 32311 32388 32404 32416
rect 32398 32376 32404 32388
rect 32456 32376 32462 32428
rect 29638 32348 29644 32360
rect 28368 32320 29224 32348
rect 29599 32320 29644 32348
rect 25240 32252 27844 32280
rect 27893 32283 27951 32289
rect 12768 32184 12848 32212
rect 12768 32172 12774 32184
rect 13906 32172 13912 32224
rect 13964 32212 13970 32224
rect 15565 32215 15623 32221
rect 15565 32212 15577 32215
rect 13964 32184 15577 32212
rect 13964 32172 13970 32184
rect 15565 32181 15577 32184
rect 15611 32181 15623 32215
rect 15565 32175 15623 32181
rect 22922 32172 22928 32224
rect 22980 32212 22986 32224
rect 23201 32215 23259 32221
rect 23201 32212 23213 32215
rect 22980 32184 23213 32212
rect 22980 32172 22986 32184
rect 23201 32181 23213 32184
rect 23247 32212 23259 32215
rect 25240 32212 25268 32252
rect 27893 32249 27905 32283
rect 27939 32280 27951 32283
rect 28902 32280 28908 32292
rect 27939 32252 28908 32280
rect 27939 32249 27951 32252
rect 27893 32243 27951 32249
rect 28902 32240 28908 32252
rect 28960 32240 28966 32292
rect 29196 32289 29224 32320
rect 29638 32308 29644 32320
rect 29696 32308 29702 32360
rect 29822 32348 29828 32360
rect 29783 32320 29828 32348
rect 29822 32308 29828 32320
rect 29880 32308 29886 32360
rect 30098 32308 30104 32360
rect 30156 32348 30162 32360
rect 32416 32348 32444 32376
rect 30156 32320 32444 32348
rect 30156 32308 30162 32320
rect 29181 32283 29239 32289
rect 29181 32249 29193 32283
rect 29227 32249 29239 32283
rect 29181 32243 29239 32249
rect 30653 32283 30711 32289
rect 30653 32249 30665 32283
rect 30699 32280 30711 32283
rect 31754 32280 31760 32292
rect 30699 32252 31760 32280
rect 30699 32249 30711 32252
rect 30653 32243 30711 32249
rect 31754 32240 31760 32252
rect 31812 32240 31818 32292
rect 23247 32184 25268 32212
rect 23247 32181 23259 32184
rect 23201 32175 23259 32181
rect 25314 32172 25320 32224
rect 25372 32212 25378 32224
rect 25869 32215 25927 32221
rect 25869 32212 25881 32215
rect 25372 32184 25881 32212
rect 25372 32172 25378 32184
rect 25869 32181 25881 32184
rect 25915 32212 25927 32215
rect 26142 32212 26148 32224
rect 25915 32184 26148 32212
rect 25915 32181 25927 32184
rect 25869 32175 25927 32181
rect 26142 32172 26148 32184
rect 26200 32172 26206 32224
rect 26786 32172 26792 32224
rect 26844 32212 26850 32224
rect 28626 32212 28632 32224
rect 26844 32184 28632 32212
rect 26844 32172 26850 32184
rect 28626 32172 28632 32184
rect 28684 32172 28690 32224
rect 28721 32215 28779 32221
rect 28721 32181 28733 32215
rect 28767 32212 28779 32215
rect 30190 32212 30196 32224
rect 28767 32184 30196 32212
rect 28767 32181 28779 32184
rect 28721 32175 28779 32181
rect 30190 32172 30196 32184
rect 30248 32172 30254 32224
rect 32585 32215 32643 32221
rect 32585 32181 32597 32215
rect 32631 32212 32643 32215
rect 32766 32212 32772 32224
rect 32631 32184 32772 32212
rect 32631 32181 32643 32184
rect 32585 32175 32643 32181
rect 32766 32172 32772 32184
rect 32824 32172 32830 32224
rect 1104 32122 48852 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 48852 32122
rect 1104 32048 48852 32070
rect 4062 31968 4068 32020
rect 4120 32008 4126 32020
rect 10870 32008 10876 32020
rect 4120 31980 10548 32008
rect 10831 31980 10876 32008
rect 4120 31968 4126 31980
rect 2958 31940 2964 31952
rect 1412 31912 2964 31940
rect 1412 31881 1440 31912
rect 2958 31900 2964 31912
rect 3016 31900 3022 31952
rect 10520 31940 10548 31980
rect 10870 31968 10876 31980
rect 10928 31968 10934 32020
rect 21910 32008 21916 32020
rect 10980 31980 17264 32008
rect 21871 31980 21916 32008
rect 10980 31940 11008 31980
rect 10520 31912 11008 31940
rect 11238 31900 11244 31952
rect 11296 31900 11302 31952
rect 13170 31900 13176 31952
rect 13228 31940 13234 31952
rect 13541 31943 13599 31949
rect 13541 31940 13553 31943
rect 13228 31912 13553 31940
rect 13228 31900 13234 31912
rect 13541 31909 13553 31912
rect 13587 31940 13599 31943
rect 17236 31940 17264 31980
rect 21910 31968 21916 31980
rect 21968 31968 21974 32020
rect 22250 31980 24992 32008
rect 22250 31940 22278 31980
rect 13587 31912 14136 31940
rect 17236 31912 22278 31940
rect 24964 31940 24992 31980
rect 25682 31968 25688 32020
rect 25740 32008 25746 32020
rect 25740 31980 28212 32008
rect 25740 31968 25746 31980
rect 27617 31943 27675 31949
rect 27617 31940 27629 31943
rect 24964 31912 26464 31940
rect 13587 31909 13599 31912
rect 13541 31903 13599 31909
rect 1397 31875 1455 31881
rect 1397 31841 1409 31875
rect 1443 31841 1455 31875
rect 1397 31835 1455 31841
rect 1581 31875 1639 31881
rect 1581 31841 1593 31875
rect 1627 31872 1639 31875
rect 3881 31875 3939 31881
rect 3881 31872 3893 31875
rect 1627 31844 3893 31872
rect 1627 31841 1639 31844
rect 1581 31835 1639 31841
rect 3881 31841 3893 31844
rect 3927 31841 3939 31875
rect 10134 31872 10140 31884
rect 10095 31844 10140 31872
rect 3881 31835 3939 31841
rect 10134 31832 10140 31844
rect 10192 31832 10198 31884
rect 3234 31804 3240 31816
rect 3195 31776 3240 31804
rect 3234 31764 3240 31776
rect 3292 31764 3298 31816
rect 3786 31804 3792 31816
rect 3747 31776 3792 31804
rect 3786 31764 3792 31776
rect 3844 31764 3850 31816
rect 10045 31807 10103 31813
rect 10045 31773 10057 31807
rect 10091 31804 10103 31807
rect 10870 31804 10876 31816
rect 10091 31776 10876 31804
rect 10091 31773 10103 31776
rect 10045 31767 10103 31773
rect 10870 31764 10876 31776
rect 10928 31764 10934 31816
rect 11146 31804 11152 31816
rect 11107 31776 11152 31804
rect 11146 31764 11152 31776
rect 11204 31764 11210 31816
rect 11253 31813 11281 31900
rect 14108 31881 14136 31912
rect 14093 31875 14151 31881
rect 14093 31841 14105 31875
rect 14139 31841 14151 31875
rect 14366 31872 14372 31884
rect 14327 31844 14372 31872
rect 14093 31835 14151 31841
rect 14366 31832 14372 31844
rect 14424 31832 14430 31884
rect 17954 31872 17960 31884
rect 17052 31844 17960 31872
rect 11238 31807 11296 31813
rect 11238 31773 11250 31807
rect 11284 31773 11296 31807
rect 11238 31767 11296 31773
rect 11333 31807 11391 31813
rect 11333 31773 11345 31807
rect 11379 31773 11391 31807
rect 11333 31767 11391 31773
rect 11348 31736 11376 31767
rect 11514 31764 11520 31816
rect 11572 31804 11578 31816
rect 12161 31807 12219 31813
rect 11572 31776 12112 31804
rect 11572 31764 11578 31776
rect 10428 31708 11376 31736
rect 10428 31677 10456 31708
rect 10413 31671 10471 31677
rect 10413 31637 10425 31671
rect 10459 31637 10471 31671
rect 12084 31668 12112 31776
rect 12161 31773 12173 31807
rect 12207 31804 12219 31807
rect 12710 31804 12716 31816
rect 12207 31776 12716 31804
rect 12207 31773 12219 31776
rect 12161 31767 12219 31773
rect 12710 31764 12716 31776
rect 12768 31764 12774 31816
rect 17052 31813 17080 31844
rect 17954 31832 17960 31844
rect 18012 31832 18018 31884
rect 19334 31832 19340 31884
rect 19392 31832 19398 31884
rect 20254 31832 20260 31884
rect 20312 31872 20318 31884
rect 21082 31872 21088 31884
rect 20312 31844 21088 31872
rect 20312 31832 20318 31844
rect 21082 31832 21088 31844
rect 21140 31832 21146 31884
rect 22646 31872 22652 31884
rect 22066 31844 22652 31872
rect 17037 31807 17095 31813
rect 17037 31773 17049 31807
rect 17083 31773 17095 31807
rect 17218 31804 17224 31816
rect 17179 31776 17224 31804
rect 17037 31767 17095 31773
rect 17218 31764 17224 31776
rect 17276 31764 17282 31816
rect 17681 31807 17739 31813
rect 17681 31773 17693 31807
rect 17727 31804 17739 31807
rect 17862 31804 17868 31816
rect 17727 31776 17761 31804
rect 17823 31776 17868 31804
rect 17727 31773 17739 31776
rect 17681 31767 17739 31773
rect 12428 31739 12486 31745
rect 12428 31705 12440 31739
rect 12474 31736 12486 31739
rect 13078 31736 13084 31748
rect 12474 31708 13084 31736
rect 12474 31705 12486 31708
rect 12428 31699 12486 31705
rect 13078 31696 13084 31708
rect 13136 31696 13142 31748
rect 17696 31736 17724 31767
rect 17862 31764 17868 31776
rect 17920 31764 17926 31816
rect 18049 31807 18107 31813
rect 18049 31773 18061 31807
rect 18095 31804 18107 31807
rect 19352 31804 19380 31832
rect 20625 31807 20683 31813
rect 20625 31804 20637 31807
rect 18095 31776 20637 31804
rect 18095 31773 18107 31776
rect 18049 31767 18107 31773
rect 20625 31773 20637 31776
rect 20671 31773 20683 31807
rect 20625 31767 20683 31773
rect 20901 31807 20959 31813
rect 20901 31773 20913 31807
rect 20947 31804 20959 31807
rect 20990 31804 20996 31816
rect 20947 31776 20996 31804
rect 20947 31773 20959 31776
rect 20901 31767 20959 31773
rect 20990 31764 20996 31776
rect 21048 31764 21054 31816
rect 22066 31804 22094 31844
rect 22646 31832 22652 31844
rect 22704 31832 22710 31884
rect 26145 31875 26203 31881
rect 26145 31841 26157 31875
rect 26191 31872 26203 31875
rect 26326 31872 26332 31884
rect 26191 31844 26332 31872
rect 26191 31841 26203 31844
rect 26145 31835 26203 31841
rect 26326 31832 26332 31844
rect 26384 31832 26390 31884
rect 22143 31807 22201 31813
rect 22143 31804 22155 31807
rect 22066 31776 22155 31804
rect 22143 31773 22155 31776
rect 22189 31773 22201 31807
rect 22143 31767 22201 31773
rect 22262 31804 22320 31810
rect 22370 31807 22376 31816
rect 22262 31770 22274 31804
rect 22308 31770 22320 31804
rect 22262 31764 22320 31770
rect 22362 31801 22376 31807
rect 22362 31767 22374 31801
rect 22362 31764 22376 31767
rect 22428 31764 22434 31816
rect 22557 31807 22615 31813
rect 22557 31773 22569 31807
rect 22603 31804 22615 31807
rect 23474 31804 23480 31816
rect 22603 31776 23480 31804
rect 22603 31773 22615 31776
rect 22557 31767 22615 31773
rect 23474 31764 23480 31776
rect 23532 31764 23538 31816
rect 25222 31764 25228 31816
rect 25280 31804 25286 31816
rect 26234 31804 26240 31816
rect 25280 31776 26240 31804
rect 25280 31764 25286 31776
rect 26234 31764 26240 31776
rect 26292 31764 26298 31816
rect 26436 31813 26464 31912
rect 26712 31912 27629 31940
rect 26421 31807 26479 31813
rect 26421 31773 26433 31807
rect 26467 31773 26479 31807
rect 26421 31767 26479 31773
rect 26513 31807 26571 31813
rect 26513 31773 26525 31807
rect 26559 31773 26571 31807
rect 26513 31767 26571 31773
rect 26626 31807 26684 31813
rect 26626 31773 26638 31807
rect 26672 31804 26684 31807
rect 26712 31804 26740 31912
rect 27617 31909 27629 31912
rect 27663 31909 27675 31943
rect 27617 31903 27675 31909
rect 27154 31832 27160 31884
rect 27212 31872 27218 31884
rect 28184 31872 28212 31980
rect 28350 31968 28356 32020
rect 28408 32008 28414 32020
rect 29730 32008 29736 32020
rect 28408 31980 29736 32008
rect 28408 31968 28414 31980
rect 29730 31968 29736 31980
rect 29788 31968 29794 32020
rect 31757 32011 31815 32017
rect 31757 31977 31769 32011
rect 31803 32008 31815 32011
rect 31846 32008 31852 32020
rect 31803 31980 31852 32008
rect 31803 31977 31815 31980
rect 31757 31971 31815 31977
rect 31846 31968 31852 31980
rect 31904 31968 31910 32020
rect 33870 32008 33876 32020
rect 33831 31980 33876 32008
rect 33870 31968 33876 31980
rect 33928 32008 33934 32020
rect 34330 32008 34336 32020
rect 33928 31980 34336 32008
rect 33928 31968 33934 31980
rect 34330 31968 34336 31980
rect 34388 31968 34394 32020
rect 35342 32008 35348 32020
rect 35303 31980 35348 32008
rect 35342 31968 35348 31980
rect 35400 31968 35406 32020
rect 28537 31875 28595 31881
rect 28537 31872 28549 31875
rect 27212 31844 27660 31872
rect 28184 31844 28549 31872
rect 27212 31832 27218 31844
rect 26672 31776 26740 31804
rect 26672 31773 26684 31776
rect 26626 31767 26684 31773
rect 17954 31736 17960 31748
rect 17696 31708 17960 31736
rect 17954 31696 17960 31708
rect 18012 31696 18018 31748
rect 19426 31696 19432 31748
rect 19484 31736 19490 31748
rect 22002 31736 22008 31748
rect 19484 31708 22008 31736
rect 19484 31696 19490 31708
rect 22002 31696 22008 31708
rect 22060 31736 22066 31748
rect 22277 31736 22305 31764
rect 22362 31761 22420 31764
rect 22060 31708 22305 31736
rect 22060 31696 22066 31708
rect 25130 31696 25136 31748
rect 25188 31736 25194 31748
rect 26528 31736 26556 31767
rect 26786 31764 26792 31816
rect 26844 31804 26850 31816
rect 27632 31804 27660 31844
rect 28537 31841 28549 31844
rect 28583 31841 28595 31875
rect 28537 31835 28595 31841
rect 28721 31875 28779 31881
rect 28721 31841 28733 31875
rect 28767 31872 28779 31875
rect 28902 31872 28908 31884
rect 28767 31844 28908 31872
rect 28767 31841 28779 31844
rect 28721 31835 28779 31841
rect 28902 31832 28908 31844
rect 28960 31872 28966 31884
rect 29822 31872 29828 31884
rect 28960 31844 29828 31872
rect 28960 31832 28966 31844
rect 29822 31832 29828 31844
rect 29880 31832 29886 31884
rect 30377 31875 30435 31881
rect 30377 31841 30389 31875
rect 30423 31841 30435 31875
rect 47854 31872 47860 31884
rect 47815 31844 47860 31872
rect 30377 31835 30435 31841
rect 30392 31804 30420 31835
rect 47854 31832 47860 31844
rect 47912 31832 47918 31884
rect 26844 31776 26889 31804
rect 27632 31801 27936 31804
rect 28184 31801 30420 31804
rect 27632 31776 30420 31801
rect 26844 31764 26850 31776
rect 27908 31773 28212 31776
rect 31754 31764 31760 31816
rect 31812 31804 31818 31816
rect 32493 31807 32551 31813
rect 32493 31804 32505 31807
rect 31812 31776 32505 31804
rect 31812 31764 31818 31776
rect 32493 31773 32505 31776
rect 32539 31773 32551 31807
rect 32493 31767 32551 31773
rect 35253 31807 35311 31813
rect 35253 31773 35265 31807
rect 35299 31804 35311 31807
rect 37274 31804 37280 31816
rect 35299 31776 37280 31804
rect 35299 31773 35311 31776
rect 35253 31767 35311 31773
rect 37274 31764 37280 31776
rect 37332 31764 37338 31816
rect 47486 31804 47492 31816
rect 47447 31776 47492 31804
rect 47486 31764 47492 31776
rect 47544 31764 47550 31816
rect 25188 31708 26556 31736
rect 27249 31739 27307 31745
rect 25188 31696 25194 31708
rect 27249 31705 27261 31739
rect 27295 31705 27307 31739
rect 27249 31699 27307 31705
rect 27433 31739 27491 31745
rect 27433 31705 27445 31739
rect 27479 31736 27491 31739
rect 28350 31736 28356 31748
rect 27479 31708 28356 31736
rect 27479 31705 27491 31708
rect 27433 31699 27491 31705
rect 14734 31668 14740 31680
rect 12084 31640 14740 31668
rect 10413 31631 10471 31637
rect 14734 31628 14740 31640
rect 14792 31668 14798 31680
rect 22462 31668 22468 31680
rect 14792 31640 22468 31668
rect 14792 31628 14798 31640
rect 22462 31628 22468 31640
rect 22520 31628 22526 31680
rect 25774 31628 25780 31680
rect 25832 31668 25838 31680
rect 27154 31668 27160 31680
rect 25832 31640 27160 31668
rect 25832 31628 25838 31640
rect 27154 31628 27160 31640
rect 27212 31628 27218 31680
rect 27264 31668 27292 31699
rect 28350 31696 28356 31708
rect 28408 31696 28414 31748
rect 29546 31736 29552 31748
rect 29507 31708 29552 31736
rect 29546 31696 29552 31708
rect 29604 31696 29610 31748
rect 29730 31736 29736 31748
rect 29691 31708 29736 31736
rect 29730 31696 29736 31708
rect 29788 31696 29794 31748
rect 30466 31696 30472 31748
rect 30524 31736 30530 31748
rect 30622 31739 30680 31745
rect 30622 31736 30634 31739
rect 30524 31708 30634 31736
rect 30524 31696 30530 31708
rect 30622 31705 30634 31708
rect 30668 31705 30680 31739
rect 30622 31699 30680 31705
rect 32122 31696 32128 31748
rect 32180 31736 32186 31748
rect 32738 31739 32796 31745
rect 32738 31736 32750 31739
rect 32180 31708 32750 31736
rect 32180 31696 32186 31708
rect 32738 31705 32750 31708
rect 32784 31705 32796 31739
rect 32738 31699 32796 31705
rect 28077 31671 28135 31677
rect 28077 31668 28089 31671
rect 27264 31640 28089 31668
rect 28077 31637 28089 31640
rect 28123 31637 28135 31671
rect 28077 31631 28135 31637
rect 28445 31671 28503 31677
rect 28445 31637 28457 31671
rect 28491 31668 28503 31671
rect 29086 31668 29092 31680
rect 28491 31640 29092 31668
rect 28491 31637 28503 31640
rect 28445 31631 28503 31637
rect 29086 31628 29092 31640
rect 29144 31628 29150 31680
rect 29917 31671 29975 31677
rect 29917 31637 29929 31671
rect 29963 31668 29975 31671
rect 30006 31668 30012 31680
rect 29963 31640 30012 31668
rect 29963 31637 29975 31640
rect 29917 31631 29975 31637
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 1104 31578 48852 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 48852 31578
rect 1104 31504 48852 31526
rect 13078 31464 13084 31476
rect 13039 31436 13084 31464
rect 13078 31424 13084 31436
rect 13136 31424 13142 31476
rect 13262 31424 13268 31476
rect 13320 31464 13326 31476
rect 13449 31467 13507 31473
rect 13449 31464 13461 31467
rect 13320 31436 13461 31464
rect 13320 31424 13326 31436
rect 13449 31433 13461 31436
rect 13495 31433 13507 31467
rect 13449 31427 13507 31433
rect 13541 31467 13599 31473
rect 13541 31433 13553 31467
rect 13587 31464 13599 31467
rect 13587 31436 13676 31464
rect 13587 31433 13599 31436
rect 13541 31427 13599 31433
rect 1486 31396 1492 31408
rect 1447 31368 1492 31396
rect 1486 31356 1492 31368
rect 1544 31356 1550 31408
rect 2317 31399 2375 31405
rect 2317 31365 2329 31399
rect 2363 31396 2375 31399
rect 3050 31396 3056 31408
rect 2363 31368 3056 31396
rect 2363 31365 2375 31368
rect 2317 31359 2375 31365
rect 3050 31356 3056 31368
rect 3108 31356 3114 31408
rect 5258 31356 5264 31408
rect 5316 31396 5322 31408
rect 12986 31396 12992 31408
rect 5316 31368 12992 31396
rect 5316 31356 5322 31368
rect 12986 31356 12992 31368
rect 13044 31356 13050 31408
rect 13648 31396 13676 31436
rect 14090 31424 14096 31476
rect 14148 31464 14154 31476
rect 14148 31436 20760 31464
rect 14148 31424 14154 31436
rect 14645 31399 14703 31405
rect 14645 31396 14657 31399
rect 13648 31368 14657 31396
rect 14645 31365 14657 31368
rect 14691 31365 14703 31399
rect 14645 31359 14703 31365
rect 14734 31356 14740 31408
rect 14792 31396 14798 31408
rect 20254 31396 20260 31408
rect 14792 31368 20260 31396
rect 14792 31356 14798 31368
rect 20254 31356 20260 31368
rect 20312 31356 20318 31408
rect 20349 31399 20407 31405
rect 20349 31365 20361 31399
rect 20395 31396 20407 31399
rect 20622 31396 20628 31408
rect 20395 31368 20628 31396
rect 20395 31365 20407 31368
rect 20349 31359 20407 31365
rect 20622 31356 20628 31368
rect 20680 31356 20686 31408
rect 20732 31396 20760 31436
rect 20990 31424 20996 31476
rect 21048 31464 21054 31476
rect 22281 31467 22339 31473
rect 21048 31436 21772 31464
rect 21048 31424 21054 31436
rect 20732 31368 21677 31396
rect 13354 31328 13360 31340
rect 13315 31300 13360 31328
rect 13354 31288 13360 31300
rect 13412 31288 13418 31340
rect 13464 31300 13952 31328
rect 2133 31263 2191 31269
rect 2133 31229 2145 31263
rect 2179 31229 2191 31263
rect 3142 31260 3148 31272
rect 3103 31232 3148 31260
rect 2133 31223 2191 31229
rect 2148 31192 2176 31223
rect 3142 31220 3148 31232
rect 3200 31220 3206 31272
rect 13464 31260 13492 31300
rect 13814 31260 13820 31272
rect 12406 31232 13492 31260
rect 13775 31232 13820 31260
rect 2866 31192 2872 31204
rect 2148 31164 2872 31192
rect 2866 31152 2872 31164
rect 2924 31152 2930 31204
rect 1581 31127 1639 31133
rect 1581 31093 1593 31127
rect 1627 31124 1639 31127
rect 12406 31124 12434 31232
rect 13814 31220 13820 31232
rect 13872 31220 13878 31272
rect 13924 31260 13952 31300
rect 13998 31288 14004 31340
rect 14056 31328 14062 31340
rect 14277 31331 14335 31337
rect 14277 31328 14289 31331
rect 14056 31300 14289 31328
rect 14056 31288 14062 31300
rect 14277 31297 14289 31300
rect 14323 31297 14335 31331
rect 14277 31291 14335 31297
rect 14366 31288 14372 31340
rect 14424 31328 14430 31340
rect 14461 31331 14519 31337
rect 14461 31328 14473 31331
rect 14424 31300 14473 31328
rect 14424 31288 14430 31300
rect 14461 31297 14473 31300
rect 14507 31297 14519 31331
rect 14461 31291 14519 31297
rect 16758 31288 16764 31340
rect 16816 31328 16822 31340
rect 16925 31331 16983 31337
rect 16925 31328 16937 31331
rect 16816 31300 16937 31328
rect 16816 31288 16822 31300
rect 16925 31297 16937 31300
rect 16971 31297 16983 31331
rect 16925 31291 16983 31297
rect 18782 31288 18788 31340
rect 18840 31328 18846 31340
rect 19242 31328 19248 31340
rect 18840 31300 19248 31328
rect 18840 31288 18846 31300
rect 19242 31288 19248 31300
rect 19300 31328 19306 31340
rect 19705 31331 19763 31337
rect 19705 31328 19717 31331
rect 19300 31300 19717 31328
rect 19300 31288 19306 31300
rect 19705 31297 19717 31300
rect 19751 31297 19763 31331
rect 19705 31291 19763 31297
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31328 20591 31331
rect 20990 31328 20996 31340
rect 20579 31300 20996 31328
rect 20579 31297 20591 31300
rect 20533 31291 20591 31297
rect 20990 31288 20996 31300
rect 21048 31288 21054 31340
rect 15102 31260 15108 31272
rect 13924 31232 15108 31260
rect 15102 31220 15108 31232
rect 15160 31220 15166 31272
rect 15194 31220 15200 31272
rect 15252 31260 15258 31272
rect 16669 31263 16727 31269
rect 16669 31260 16681 31263
rect 15252 31232 16681 31260
rect 15252 31220 15258 31232
rect 16669 31229 16681 31232
rect 16715 31229 16727 31263
rect 16669 31223 16727 31229
rect 20717 31263 20775 31269
rect 20717 31229 20729 31263
rect 20763 31260 20775 31263
rect 20806 31260 20812 31272
rect 20763 31232 20812 31260
rect 20763 31229 20775 31232
rect 20717 31223 20775 31229
rect 20806 31220 20812 31232
rect 20864 31220 20870 31272
rect 21649 31260 21677 31368
rect 21744 31328 21772 31436
rect 22281 31433 22293 31467
rect 22327 31464 22339 31467
rect 22370 31464 22376 31476
rect 22327 31436 22376 31464
rect 22327 31433 22339 31436
rect 22281 31427 22339 31433
rect 22370 31424 22376 31436
rect 22428 31424 22434 31476
rect 22462 31424 22468 31476
rect 22520 31464 22526 31476
rect 24302 31464 24308 31476
rect 22520 31436 24164 31464
rect 24263 31436 24308 31464
rect 22520 31424 22526 31436
rect 21913 31399 21971 31405
rect 21913 31365 21925 31399
rect 21959 31396 21971 31399
rect 22186 31396 22192 31408
rect 21959 31368 22192 31396
rect 21959 31365 21971 31368
rect 21913 31359 21971 31365
rect 22186 31356 22192 31368
rect 22244 31356 22250 31408
rect 23201 31399 23259 31405
rect 23201 31396 23213 31399
rect 22296 31368 23213 31396
rect 22097 31331 22155 31337
rect 22097 31328 22109 31331
rect 21744 31300 22109 31328
rect 22097 31297 22109 31300
rect 22143 31328 22155 31331
rect 22296 31328 22324 31368
rect 23201 31365 23213 31368
rect 23247 31396 23259 31399
rect 23290 31396 23296 31408
rect 23247 31368 23296 31396
rect 23247 31365 23259 31368
rect 23201 31359 23259 31365
rect 23290 31356 23296 31368
rect 23348 31356 23354 31408
rect 24136 31396 24164 31436
rect 24302 31424 24308 31436
rect 24360 31424 24366 31476
rect 25225 31467 25283 31473
rect 25225 31433 25237 31467
rect 25271 31464 25283 31467
rect 26786 31464 26792 31476
rect 25271 31436 26792 31464
rect 25271 31433 25283 31436
rect 25225 31427 25283 31433
rect 26786 31424 26792 31436
rect 26844 31424 26850 31476
rect 28537 31467 28595 31473
rect 28537 31433 28549 31467
rect 28583 31464 28595 31467
rect 29546 31464 29552 31476
rect 28583 31436 29552 31464
rect 28583 31433 28595 31436
rect 28537 31427 28595 31433
rect 29546 31424 29552 31436
rect 29604 31424 29610 31476
rect 29733 31467 29791 31473
rect 29733 31433 29745 31467
rect 29779 31464 29791 31467
rect 30466 31464 30472 31476
rect 29779 31436 30472 31464
rect 29779 31433 29791 31436
rect 29733 31427 29791 31433
rect 30466 31424 30472 31436
rect 30524 31424 30530 31476
rect 32122 31464 32128 31476
rect 32083 31436 32128 31464
rect 32122 31424 32128 31436
rect 32180 31424 32186 31476
rect 24762 31396 24768 31408
rect 24136 31368 24768 31396
rect 24762 31356 24768 31368
rect 24820 31356 24826 31408
rect 26234 31356 26240 31408
rect 26292 31396 26298 31408
rect 26418 31396 26424 31408
rect 26292 31368 26424 31396
rect 26292 31356 26298 31368
rect 26418 31356 26424 31368
rect 26476 31356 26482 31408
rect 27065 31399 27123 31405
rect 27065 31365 27077 31399
rect 27111 31396 27123 31399
rect 27890 31396 27896 31408
rect 27111 31368 27896 31396
rect 27111 31365 27123 31368
rect 27065 31359 27123 31365
rect 27890 31356 27896 31368
rect 27948 31356 27954 31408
rect 28810 31356 28816 31408
rect 28868 31396 28874 31408
rect 28868 31368 30604 31396
rect 28868 31356 28874 31368
rect 23014 31328 23020 31340
rect 22143 31300 22324 31328
rect 22975 31300 23020 31328
rect 22143 31297 22155 31300
rect 22097 31291 22155 31297
rect 23014 31288 23020 31300
rect 23072 31288 23078 31340
rect 24026 31288 24032 31340
rect 24084 31328 24090 31340
rect 24213 31331 24271 31337
rect 24213 31328 24225 31331
rect 24084 31300 24225 31328
rect 24084 31288 24090 31300
rect 24213 31297 24225 31300
rect 24259 31328 24271 31331
rect 24394 31328 24400 31340
rect 24259 31300 24400 31328
rect 24259 31297 24271 31300
rect 24213 31291 24271 31297
rect 24394 31288 24400 31300
rect 24452 31288 24458 31340
rect 25133 31331 25191 31337
rect 25133 31297 25145 31331
rect 25179 31297 25191 31331
rect 25133 31291 25191 31297
rect 25869 31331 25927 31337
rect 25869 31297 25881 31331
rect 25915 31297 25927 31331
rect 25869 31291 25927 31297
rect 28905 31331 28963 31337
rect 28905 31297 28917 31331
rect 28951 31328 28963 31331
rect 29638 31328 29644 31340
rect 28951 31300 29644 31328
rect 28951 31297 28963 31300
rect 28905 31291 28963 31297
rect 23106 31260 23112 31272
rect 21649 31232 23112 31260
rect 23106 31220 23112 31232
rect 23164 31220 23170 31272
rect 23842 31220 23848 31272
rect 23900 31260 23906 31272
rect 25038 31260 25044 31272
rect 23900 31232 25044 31260
rect 23900 31220 23906 31232
rect 25038 31220 25044 31232
rect 25096 31260 25102 31272
rect 25148 31260 25176 31291
rect 25096 31232 25176 31260
rect 25096 31220 25102 31232
rect 12710 31152 12716 31204
rect 12768 31192 12774 31204
rect 15212 31192 15240 31220
rect 12768 31164 15240 31192
rect 19889 31195 19947 31201
rect 12768 31152 12774 31164
rect 19889 31161 19901 31195
rect 19935 31192 19947 31195
rect 20162 31192 20168 31204
rect 19935 31164 20168 31192
rect 19935 31161 19947 31164
rect 19889 31155 19947 31161
rect 20162 31152 20168 31164
rect 20220 31192 20226 31204
rect 21358 31192 21364 31204
rect 20220 31164 21364 31192
rect 20220 31152 20226 31164
rect 21358 31152 21364 31164
rect 21416 31152 21422 31204
rect 25884 31192 25912 31291
rect 29638 31288 29644 31300
rect 29696 31288 29702 31340
rect 30009 31331 30067 31337
rect 30009 31328 30021 31331
rect 29840 31300 30021 31328
rect 26142 31220 26148 31272
rect 26200 31260 26206 31272
rect 28997 31263 29055 31269
rect 28997 31260 29009 31263
rect 26200 31232 29009 31260
rect 26200 31220 26206 31232
rect 28997 31229 29009 31232
rect 29043 31229 29055 31263
rect 28997 31223 29055 31229
rect 29089 31263 29147 31269
rect 29089 31229 29101 31263
rect 29135 31229 29147 31263
rect 29089 31223 29147 31229
rect 23216 31164 25912 31192
rect 25976 31164 28856 31192
rect 13722 31124 13728 31136
rect 1627 31096 12434 31124
rect 13635 31096 13728 31124
rect 1627 31093 1639 31096
rect 1581 31087 1639 31093
rect 13722 31084 13728 31096
rect 13780 31124 13786 31136
rect 14458 31124 14464 31136
rect 13780 31096 14464 31124
rect 13780 31084 13786 31096
rect 14458 31084 14464 31096
rect 14516 31084 14522 31136
rect 18046 31124 18052 31136
rect 18007 31096 18052 31124
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 19242 31084 19248 31136
rect 19300 31124 19306 31136
rect 23216 31124 23244 31164
rect 25976 31136 26004 31164
rect 19300 31096 23244 31124
rect 19300 31084 19306 31096
rect 23290 31084 23296 31136
rect 23348 31124 23354 31136
rect 23385 31127 23443 31133
rect 23385 31124 23397 31127
rect 23348 31096 23397 31124
rect 23348 31084 23354 31096
rect 23385 31093 23397 31096
rect 23431 31093 23443 31127
rect 25958 31124 25964 31136
rect 25919 31096 25964 31124
rect 23385 31087 23443 31093
rect 25958 31084 25964 31096
rect 26016 31084 26022 31136
rect 26970 31084 26976 31136
rect 27028 31124 27034 31136
rect 27154 31124 27160 31136
rect 27028 31096 27160 31124
rect 27028 31084 27034 31096
rect 27154 31084 27160 31096
rect 27212 31084 27218 31136
rect 28828 31124 28856 31164
rect 28902 31152 28908 31204
rect 28960 31192 28966 31204
rect 29104 31192 29132 31223
rect 29730 31220 29736 31272
rect 29788 31260 29794 31272
rect 29840 31260 29868 31300
rect 30009 31297 30021 31300
rect 30055 31297 30067 31331
rect 30009 31291 30067 31297
rect 30101 31331 30159 31337
rect 30101 31297 30113 31331
rect 30147 31297 30159 31331
rect 30101 31291 30159 31297
rect 30116 31260 30144 31291
rect 30190 31288 30196 31340
rect 30248 31328 30254 31340
rect 30248 31300 30293 31328
rect 30248 31288 30254 31300
rect 30374 31288 30380 31340
rect 30432 31328 30438 31340
rect 30432 31300 30477 31328
rect 30432 31288 30438 31300
rect 29788 31232 29868 31260
rect 30024 31232 30144 31260
rect 30576 31260 30604 31368
rect 31846 31356 31852 31408
rect 31904 31396 31910 31408
rect 31904 31368 32536 31396
rect 31904 31356 31910 31368
rect 30926 31288 30932 31340
rect 30984 31328 30990 31340
rect 32508 31337 32536 31368
rect 32401 31331 32459 31337
rect 32401 31328 32413 31331
rect 30984 31300 32413 31328
rect 30984 31288 30990 31300
rect 32401 31297 32413 31300
rect 32447 31297 32459 31331
rect 32401 31291 32459 31297
rect 32493 31331 32551 31337
rect 32493 31297 32505 31331
rect 32539 31297 32551 31331
rect 32493 31291 32551 31297
rect 32582 31288 32588 31340
rect 32640 31328 32646 31340
rect 32766 31328 32772 31340
rect 32640 31300 32685 31328
rect 32727 31300 32772 31328
rect 32640 31288 32646 31300
rect 32766 31288 32772 31300
rect 32824 31288 32830 31340
rect 47946 31328 47952 31340
rect 47907 31300 47952 31328
rect 47946 31288 47952 31300
rect 48004 31288 48010 31340
rect 48133 31263 48191 31269
rect 48133 31260 48145 31263
rect 30576 31232 48145 31260
rect 29788 31220 29794 31232
rect 30024 31192 30052 31232
rect 48133 31229 48145 31232
rect 48179 31229 48191 31263
rect 48133 31223 48191 31229
rect 28960 31164 29132 31192
rect 29196 31164 30052 31192
rect 28960 31152 28966 31164
rect 29196 31136 29224 31164
rect 30190 31152 30196 31204
rect 30248 31192 30254 31204
rect 38838 31192 38844 31204
rect 30248 31164 38844 31192
rect 30248 31152 30254 31164
rect 38838 31152 38844 31164
rect 38896 31152 38902 31204
rect 29178 31124 29184 31136
rect 28828 31096 29184 31124
rect 29178 31084 29184 31096
rect 29236 31084 29242 31136
rect 1104 31034 48852 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 48852 31034
rect 1104 30960 48852 30982
rect 1946 30880 1952 30932
rect 2004 30920 2010 30932
rect 2317 30923 2375 30929
rect 2317 30920 2329 30923
rect 2004 30892 2329 30920
rect 2004 30880 2010 30892
rect 2317 30889 2329 30892
rect 2363 30889 2375 30923
rect 2317 30883 2375 30889
rect 2958 30880 2964 30932
rect 3016 30920 3022 30932
rect 3053 30923 3111 30929
rect 3053 30920 3065 30923
rect 3016 30892 3065 30920
rect 3016 30880 3022 30892
rect 3053 30889 3065 30892
rect 3099 30889 3111 30923
rect 3053 30883 3111 30889
rect 10134 30880 10140 30932
rect 10192 30920 10198 30932
rect 10321 30923 10379 30929
rect 10321 30920 10333 30923
rect 10192 30892 10333 30920
rect 10192 30880 10198 30892
rect 10321 30889 10333 30892
rect 10367 30889 10379 30923
rect 16850 30920 16856 30932
rect 16811 30892 16856 30920
rect 10321 30883 10379 30889
rect 16850 30880 16856 30892
rect 16908 30920 16914 30932
rect 17862 30920 17868 30932
rect 16908 30892 17868 30920
rect 16908 30880 16914 30892
rect 17862 30880 17868 30892
rect 17920 30880 17926 30932
rect 23014 30880 23020 30932
rect 23072 30920 23078 30932
rect 24397 30923 24455 30929
rect 24397 30920 24409 30923
rect 23072 30892 24409 30920
rect 23072 30880 23078 30892
rect 24397 30889 24409 30892
rect 24443 30889 24455 30923
rect 24397 30883 24455 30889
rect 24762 30880 24768 30932
rect 24820 30920 24826 30932
rect 24820 30892 26280 30920
rect 24820 30880 24826 30892
rect 11238 30852 11244 30864
rect 11151 30824 11244 30852
rect 11238 30812 11244 30824
rect 11296 30852 11302 30864
rect 11790 30852 11796 30864
rect 11296 30824 11796 30852
rect 11296 30812 11302 30824
rect 11790 30812 11796 30824
rect 11848 30812 11854 30864
rect 15194 30852 15200 30864
rect 15155 30824 15200 30852
rect 15194 30812 15200 30824
rect 15252 30812 15258 30864
rect 20438 30812 20444 30864
rect 20496 30852 20502 30864
rect 23474 30852 23480 30864
rect 20496 30824 23480 30852
rect 20496 30812 20502 30824
rect 2225 30719 2283 30725
rect 2225 30685 2237 30719
rect 2271 30716 2283 30719
rect 2958 30716 2964 30728
rect 2271 30688 2964 30716
rect 2271 30685 2283 30688
rect 2225 30679 2283 30685
rect 2958 30676 2964 30688
rect 3016 30676 3022 30728
rect 10042 30676 10048 30728
rect 10100 30716 10106 30728
rect 10229 30719 10287 30725
rect 10229 30716 10241 30719
rect 10100 30688 10241 30716
rect 10100 30676 10106 30688
rect 10229 30685 10241 30688
rect 10275 30685 10287 30719
rect 10410 30716 10416 30728
rect 10371 30688 10416 30716
rect 10229 30679 10287 30685
rect 10410 30676 10416 30688
rect 10468 30676 10474 30728
rect 11146 30716 11152 30728
rect 11107 30688 11152 30716
rect 11146 30676 11152 30688
rect 11204 30676 11210 30728
rect 11253 30725 11281 30812
rect 18046 30784 18052 30796
rect 16684 30756 18052 30784
rect 11238 30719 11296 30725
rect 11238 30685 11250 30719
rect 11284 30685 11296 30719
rect 11238 30679 11296 30685
rect 11333 30719 11391 30725
rect 11333 30685 11345 30719
rect 11379 30685 11391 30719
rect 11514 30716 11520 30728
rect 11475 30688 11520 30716
rect 11333 30679 11391 30685
rect 8294 30608 8300 30660
rect 8352 30648 8358 30660
rect 10873 30651 10931 30657
rect 10873 30648 10885 30651
rect 8352 30620 10885 30648
rect 8352 30608 8358 30620
rect 10873 30617 10885 30620
rect 10919 30617 10931 30651
rect 10873 30611 10931 30617
rect 9950 30540 9956 30592
rect 10008 30580 10014 30592
rect 11348 30580 11376 30679
rect 11514 30676 11520 30688
rect 11572 30676 11578 30728
rect 13906 30676 13912 30728
rect 13964 30716 13970 30728
rect 14093 30719 14151 30725
rect 14093 30716 14105 30719
rect 13964 30688 14105 30716
rect 13964 30676 13970 30688
rect 14093 30685 14105 30688
rect 14139 30685 14151 30719
rect 14274 30716 14280 30728
rect 14235 30688 14280 30716
rect 14093 30679 14151 30685
rect 14274 30676 14280 30688
rect 14332 30676 14338 30728
rect 16684 30725 16712 30756
rect 16669 30719 16727 30725
rect 16669 30685 16681 30719
rect 16715 30685 16727 30719
rect 16669 30679 16727 30685
rect 17402 30676 17408 30728
rect 17460 30716 17466 30728
rect 17788 30725 17816 30756
rect 18046 30744 18052 30756
rect 18104 30744 18110 30796
rect 20162 30744 20168 30796
rect 20220 30784 20226 30796
rect 20220 30756 20760 30784
rect 20220 30744 20226 30756
rect 20732 30725 20760 30756
rect 21008 30725 21036 30824
rect 23474 30812 23480 30824
rect 23532 30812 23538 30864
rect 24302 30812 24308 30864
rect 24360 30852 24366 30864
rect 24360 30824 24992 30852
rect 24360 30812 24366 30824
rect 21818 30744 21824 30796
rect 21876 30784 21882 30796
rect 22189 30787 22247 30793
rect 22189 30784 22201 30787
rect 21876 30756 22201 30784
rect 21876 30744 21882 30756
rect 22189 30753 22201 30756
rect 22235 30753 22247 30787
rect 24854 30784 24860 30796
rect 24815 30756 24860 30784
rect 22189 30747 22247 30753
rect 24854 30744 24860 30756
rect 24912 30744 24918 30796
rect 24964 30793 24992 30824
rect 25498 30812 25504 30864
rect 25556 30852 25562 30864
rect 25866 30852 25872 30864
rect 25556 30824 25872 30852
rect 25556 30812 25562 30824
rect 25866 30812 25872 30824
rect 25924 30812 25930 30864
rect 25958 30812 25964 30864
rect 26016 30812 26022 30864
rect 24949 30787 25007 30793
rect 24949 30753 24961 30787
rect 24995 30753 25007 30787
rect 24949 30747 25007 30753
rect 17589 30719 17647 30725
rect 17589 30716 17601 30719
rect 17460 30688 17601 30716
rect 17460 30676 17466 30688
rect 17589 30685 17601 30688
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 20579 30719 20637 30725
rect 20579 30716 20591 30719
rect 17773 30679 17831 30685
rect 20180 30688 20591 30716
rect 20180 30660 20208 30688
rect 20579 30685 20591 30688
rect 20625 30685 20637 30719
rect 20579 30679 20637 30685
rect 20714 30719 20772 30725
rect 20714 30685 20726 30719
rect 20760 30685 20772 30719
rect 20714 30679 20772 30685
rect 20809 30719 20867 30725
rect 20809 30685 20821 30719
rect 20855 30685 20867 30719
rect 20809 30679 20867 30685
rect 20993 30719 21051 30725
rect 20993 30685 21005 30719
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 22005 30719 22063 30725
rect 22005 30685 22017 30719
rect 22051 30716 22063 30719
rect 22094 30716 22100 30728
rect 22051 30688 22100 30716
rect 22051 30685 22063 30688
rect 22005 30679 22063 30685
rect 15013 30651 15071 30657
rect 15013 30617 15025 30651
rect 15059 30648 15071 30651
rect 17218 30648 17224 30660
rect 15059 30620 17224 30648
rect 15059 30617 15071 30620
rect 15013 30611 15071 30617
rect 17218 30608 17224 30620
rect 17276 30648 17282 30660
rect 19337 30651 19395 30657
rect 19337 30648 19349 30651
rect 17276 30620 19349 30648
rect 17276 30608 17282 30620
rect 19337 30617 19349 30620
rect 19383 30617 19395 30651
rect 19337 30611 19395 30617
rect 20162 30608 20168 30660
rect 20220 30608 20226 30660
rect 20824 30648 20852 30679
rect 22094 30676 22100 30688
rect 22152 30676 22158 30728
rect 23106 30716 23112 30728
rect 23067 30688 23112 30716
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 23201 30719 23259 30725
rect 23201 30685 23213 30719
rect 23247 30685 23259 30719
rect 23201 30679 23259 30685
rect 21266 30648 21272 30660
rect 20824 30620 21272 30648
rect 21266 30608 21272 30620
rect 21324 30608 21330 30660
rect 21358 30608 21364 30660
rect 21416 30648 21422 30660
rect 23216 30648 23244 30679
rect 23290 30676 23296 30728
rect 23348 30716 23354 30728
rect 23348 30688 23393 30716
rect 23348 30676 23354 30688
rect 23474 30676 23480 30728
rect 23532 30716 23538 30728
rect 23532 30688 23577 30716
rect 23532 30676 23538 30688
rect 25774 30676 25780 30728
rect 25832 30716 25838 30728
rect 25976 30725 26004 30812
rect 25869 30719 25927 30725
rect 25869 30716 25881 30719
rect 25832 30688 25881 30716
rect 25832 30676 25838 30688
rect 25869 30685 25881 30688
rect 25915 30685 25927 30719
rect 25869 30679 25927 30685
rect 25961 30719 26019 30725
rect 25961 30685 25973 30719
rect 26007 30685 26019 30719
rect 25961 30679 26019 30685
rect 26050 30676 26056 30728
rect 26108 30716 26114 30728
rect 26252 30725 26280 30892
rect 26786 30880 26792 30932
rect 26844 30920 26850 30932
rect 30190 30920 30196 30932
rect 26844 30892 30196 30920
rect 26844 30880 26850 30892
rect 30190 30880 30196 30892
rect 30248 30880 30254 30932
rect 40957 30923 41015 30929
rect 40957 30889 40969 30923
rect 41003 30920 41015 30923
rect 41506 30920 41512 30932
rect 41003 30892 41512 30920
rect 41003 30889 41015 30892
rect 40957 30883 41015 30889
rect 41506 30880 41512 30892
rect 41564 30880 41570 30932
rect 42794 30784 42800 30796
rect 29840 30756 42800 30784
rect 26237 30719 26295 30725
rect 26108 30688 26153 30716
rect 26108 30676 26114 30688
rect 26237 30685 26249 30719
rect 26283 30685 26295 30719
rect 26237 30679 26295 30685
rect 26326 30676 26332 30728
rect 26384 30716 26390 30728
rect 26970 30716 26976 30728
rect 26384 30688 26976 30716
rect 26384 30676 26390 30688
rect 26970 30676 26976 30688
rect 27028 30676 27034 30728
rect 29178 30676 29184 30728
rect 29236 30676 29242 30728
rect 29840 30725 29868 30756
rect 42794 30744 42800 30756
rect 42852 30744 42858 30796
rect 29825 30719 29883 30725
rect 29825 30685 29837 30719
rect 29871 30685 29883 30719
rect 29825 30679 29883 30685
rect 29917 30719 29975 30725
rect 29917 30685 29929 30719
rect 29963 30685 29975 30719
rect 29917 30679 29975 30685
rect 25130 30648 25136 30660
rect 21416 30620 25136 30648
rect 21416 30608 21422 30620
rect 25130 30608 25136 30620
rect 25188 30608 25194 30660
rect 26418 30608 26424 30660
rect 26476 30648 26482 30660
rect 27218 30651 27276 30657
rect 27218 30648 27230 30651
rect 26476 30620 27230 30648
rect 26476 30608 26482 30620
rect 27218 30617 27230 30620
rect 27264 30617 27276 30651
rect 29196 30648 29224 30676
rect 29932 30648 29960 30679
rect 30006 30676 30012 30728
rect 30064 30716 30070 30728
rect 30193 30719 30251 30725
rect 30064 30688 30109 30716
rect 30064 30676 30070 30688
rect 30193 30685 30205 30719
rect 30239 30716 30251 30719
rect 30282 30716 30288 30728
rect 30239 30688 30288 30716
rect 30239 30685 30251 30688
rect 30193 30679 30251 30685
rect 30282 30676 30288 30688
rect 30340 30676 30346 30728
rect 31389 30719 31447 30725
rect 31389 30685 31401 30719
rect 31435 30716 31447 30719
rect 33226 30716 33232 30728
rect 31435 30688 31754 30716
rect 33139 30688 33232 30716
rect 31435 30685 31447 30688
rect 31389 30679 31447 30685
rect 29196 30620 29960 30648
rect 31573 30651 31631 30657
rect 27218 30611 27276 30617
rect 31573 30617 31585 30651
rect 31619 30617 31631 30651
rect 31726 30648 31754 30688
rect 33226 30676 33232 30688
rect 33284 30716 33290 30728
rect 33502 30716 33508 30728
rect 33284 30688 33508 30716
rect 33284 30676 33290 30688
rect 33502 30676 33508 30688
rect 33560 30676 33566 30728
rect 33962 30716 33968 30728
rect 33923 30688 33968 30716
rect 33962 30676 33968 30688
rect 34020 30676 34026 30728
rect 34330 30676 34336 30728
rect 34388 30716 34394 30728
rect 34701 30719 34759 30725
rect 34701 30716 34713 30719
rect 34388 30688 34713 30716
rect 34388 30676 34394 30688
rect 34701 30685 34713 30688
rect 34747 30685 34759 30719
rect 34701 30679 34759 30685
rect 40126 30676 40132 30728
rect 40184 30716 40190 30728
rect 40773 30719 40831 30725
rect 40773 30716 40785 30719
rect 40184 30688 40785 30716
rect 40184 30676 40190 30688
rect 40773 30685 40785 30688
rect 40819 30685 40831 30719
rect 40773 30679 40831 30685
rect 33410 30648 33416 30660
rect 31726 30620 33416 30648
rect 31573 30611 31631 30617
rect 10008 30552 11376 30580
rect 10008 30540 10014 30552
rect 14366 30540 14372 30592
rect 14424 30580 14430 30592
rect 14461 30583 14519 30589
rect 14461 30580 14473 30583
rect 14424 30552 14473 30580
rect 14424 30540 14430 30552
rect 14461 30549 14473 30552
rect 14507 30549 14519 30583
rect 14461 30543 14519 30549
rect 16942 30540 16948 30592
rect 17000 30580 17006 30592
rect 17129 30583 17187 30589
rect 17129 30580 17141 30583
rect 17000 30552 17141 30580
rect 17000 30540 17006 30552
rect 17129 30549 17141 30552
rect 17175 30549 17187 30583
rect 17678 30580 17684 30592
rect 17639 30552 17684 30580
rect 17129 30543 17187 30549
rect 17678 30540 17684 30552
rect 17736 30540 17742 30592
rect 19426 30580 19432 30592
rect 19387 30552 19432 30580
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 20349 30583 20407 30589
rect 20349 30549 20361 30583
rect 20395 30580 20407 30583
rect 20806 30580 20812 30592
rect 20395 30552 20812 30580
rect 20395 30549 20407 30552
rect 20349 30543 20407 30549
rect 20806 30540 20812 30552
rect 20864 30540 20870 30592
rect 21634 30580 21640 30592
rect 21595 30552 21640 30580
rect 21634 30540 21640 30552
rect 21692 30540 21698 30592
rect 22097 30583 22155 30589
rect 22097 30549 22109 30583
rect 22143 30580 22155 30583
rect 22738 30580 22744 30592
rect 22143 30552 22744 30580
rect 22143 30549 22155 30552
rect 22097 30543 22155 30549
rect 22738 30540 22744 30552
rect 22796 30540 22802 30592
rect 22833 30583 22891 30589
rect 22833 30549 22845 30583
rect 22879 30580 22891 30583
rect 23014 30580 23020 30592
rect 22879 30552 23020 30580
rect 22879 30549 22891 30552
rect 22833 30543 22891 30549
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 24302 30540 24308 30592
rect 24360 30580 24366 30592
rect 24765 30583 24823 30589
rect 24765 30580 24777 30583
rect 24360 30552 24777 30580
rect 24360 30540 24366 30552
rect 24765 30549 24777 30552
rect 24811 30549 24823 30583
rect 25590 30580 25596 30592
rect 25551 30552 25596 30580
rect 24765 30543 24823 30549
rect 25590 30540 25596 30552
rect 25648 30540 25654 30592
rect 28353 30583 28411 30589
rect 28353 30549 28365 30583
rect 28399 30580 28411 30583
rect 29086 30580 29092 30592
rect 28399 30552 29092 30580
rect 28399 30549 28411 30552
rect 28353 30543 28411 30549
rect 29086 30540 29092 30552
rect 29144 30540 29150 30592
rect 29178 30540 29184 30592
rect 29236 30580 29242 30592
rect 29549 30583 29607 30589
rect 29549 30580 29561 30583
rect 29236 30552 29561 30580
rect 29236 30540 29242 30552
rect 29549 30549 29561 30552
rect 29595 30549 29607 30583
rect 31588 30580 31616 30611
rect 33410 30608 33416 30620
rect 33468 30608 33474 30660
rect 34057 30651 34115 30657
rect 34057 30617 34069 30651
rect 34103 30648 34115 30651
rect 34885 30651 34943 30657
rect 34885 30648 34897 30651
rect 34103 30620 34897 30648
rect 34103 30617 34115 30620
rect 34057 30611 34115 30617
rect 34885 30617 34897 30620
rect 34931 30617 34943 30651
rect 34885 30611 34943 30617
rect 36541 30651 36599 30657
rect 36541 30617 36553 30651
rect 36587 30648 36599 30651
rect 48498 30648 48504 30660
rect 36587 30620 48504 30648
rect 36587 30617 36599 30620
rect 36541 30611 36599 30617
rect 48498 30608 48504 30620
rect 48556 30608 48562 30660
rect 31662 30580 31668 30592
rect 31588 30552 31668 30580
rect 29549 30543 29607 30549
rect 31662 30540 31668 30552
rect 31720 30540 31726 30592
rect 31757 30583 31815 30589
rect 31757 30549 31769 30583
rect 31803 30580 31815 30583
rect 32214 30580 32220 30592
rect 31803 30552 32220 30580
rect 31803 30549 31815 30552
rect 31757 30543 31815 30549
rect 32214 30540 32220 30552
rect 32272 30540 32278 30592
rect 33321 30583 33379 30589
rect 33321 30549 33333 30583
rect 33367 30580 33379 30583
rect 33594 30580 33600 30592
rect 33367 30552 33600 30580
rect 33367 30549 33379 30552
rect 33321 30543 33379 30549
rect 33594 30540 33600 30552
rect 33652 30540 33658 30592
rect 1104 30490 48852 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 48852 30490
rect 1104 30416 48852 30438
rect 9674 30336 9680 30388
rect 9732 30376 9738 30388
rect 10410 30376 10416 30388
rect 9732 30348 10416 30376
rect 9732 30336 9738 30348
rect 10410 30336 10416 30348
rect 10468 30376 10474 30388
rect 10962 30376 10968 30388
rect 10468 30348 10968 30376
rect 10468 30336 10474 30348
rect 10962 30336 10968 30348
rect 11020 30336 11026 30388
rect 13354 30376 13360 30388
rect 13267 30348 13360 30376
rect 13354 30336 13360 30348
rect 13412 30376 13418 30388
rect 18506 30376 18512 30388
rect 13412 30348 18512 30376
rect 13412 30336 13418 30348
rect 18506 30336 18512 30348
rect 18564 30336 18570 30388
rect 21266 30376 21272 30388
rect 21227 30348 21272 30376
rect 21266 30336 21272 30348
rect 21324 30336 21330 30388
rect 23474 30336 23480 30388
rect 23532 30376 23538 30388
rect 24946 30376 24952 30388
rect 23532 30348 24952 30376
rect 23532 30336 23538 30348
rect 24946 30336 24952 30348
rect 25004 30336 25010 30388
rect 25869 30379 25927 30385
rect 25869 30345 25881 30379
rect 25915 30376 25927 30379
rect 26050 30376 26056 30388
rect 25915 30348 26056 30376
rect 25915 30345 25927 30348
rect 25869 30339 25927 30345
rect 26050 30336 26056 30348
rect 26108 30336 26114 30388
rect 29086 30336 29092 30388
rect 29144 30376 29150 30388
rect 29144 30348 31340 30376
rect 29144 30336 29150 30348
rect 8202 30308 8208 30320
rect 7760 30280 8208 30308
rect 2038 30200 2044 30252
rect 2096 30240 2102 30252
rect 7760 30249 7788 30280
rect 8202 30268 8208 30280
rect 8260 30308 8266 30320
rect 12710 30308 12716 30320
rect 8260 30280 12716 30308
rect 8260 30268 8266 30280
rect 2225 30243 2283 30249
rect 2225 30240 2237 30243
rect 2096 30212 2237 30240
rect 2096 30200 2102 30212
rect 2225 30209 2237 30212
rect 2271 30209 2283 30243
rect 2225 30203 2283 30209
rect 7745 30243 7803 30249
rect 7745 30209 7757 30243
rect 7791 30209 7803 30243
rect 7745 30203 7803 30209
rect 8012 30243 8070 30249
rect 8012 30209 8024 30243
rect 8058 30240 8070 30243
rect 8294 30240 8300 30252
rect 8058 30212 8300 30240
rect 8058 30209 8070 30212
rect 8012 30203 8070 30209
rect 8294 30200 8300 30212
rect 8352 30200 8358 30252
rect 9600 30249 9628 30280
rect 12710 30268 12716 30280
rect 12768 30268 12774 30320
rect 9585 30243 9643 30249
rect 9585 30209 9597 30243
rect 9631 30209 9643 30243
rect 9585 30203 9643 30209
rect 9852 30243 9910 30249
rect 9852 30209 9864 30243
rect 9898 30240 9910 30243
rect 10318 30240 10324 30252
rect 9898 30212 10324 30240
rect 9898 30209 9910 30212
rect 9852 30203 9910 30209
rect 10318 30200 10324 30212
rect 10376 30200 10382 30252
rect 11146 30200 11152 30252
rect 11204 30240 11210 30252
rect 13372 30249 13400 30336
rect 13449 30311 13507 30317
rect 13449 30277 13461 30311
rect 13495 30308 13507 30311
rect 14277 30311 14335 30317
rect 14277 30308 14289 30311
rect 13495 30280 14289 30308
rect 13495 30277 13507 30280
rect 13449 30271 13507 30277
rect 14277 30277 14289 30280
rect 14323 30277 14335 30311
rect 14277 30271 14335 30277
rect 14366 30268 14372 30320
rect 14424 30308 14430 30320
rect 14645 30311 14703 30317
rect 14645 30308 14657 30311
rect 14424 30280 14657 30308
rect 14424 30268 14430 30280
rect 14645 30277 14657 30280
rect 14691 30308 14703 30311
rect 15381 30311 15439 30317
rect 15381 30308 15393 30311
rect 14691 30280 15393 30308
rect 14691 30277 14703 30280
rect 14645 30271 14703 30277
rect 15381 30277 15393 30280
rect 15427 30277 15439 30311
rect 15381 30271 15439 30277
rect 16669 30311 16727 30317
rect 16669 30277 16681 30311
rect 16715 30308 16727 30311
rect 17034 30308 17040 30320
rect 16715 30280 17040 30308
rect 16715 30277 16727 30280
rect 16669 30271 16727 30277
rect 17034 30268 17040 30280
rect 17092 30268 17098 30320
rect 20901 30311 20959 30317
rect 20901 30277 20913 30311
rect 20947 30308 20959 30311
rect 21634 30308 21640 30320
rect 20947 30280 21640 30308
rect 20947 30277 20959 30280
rect 20901 30271 20959 30277
rect 21634 30268 21640 30280
rect 21692 30268 21698 30320
rect 26326 30308 26332 30320
rect 22940 30280 26332 30308
rect 13357 30243 13415 30249
rect 11204 30212 11928 30240
rect 11204 30200 11210 30212
rect 11422 30132 11428 30184
rect 11480 30172 11486 30184
rect 11900 30181 11928 30212
rect 13357 30209 13369 30243
rect 13403 30209 13415 30243
rect 13357 30203 13415 30209
rect 13541 30243 13599 30249
rect 13541 30209 13553 30243
rect 13587 30240 13599 30243
rect 14458 30240 14464 30252
rect 13587 30212 13952 30240
rect 14419 30212 14464 30240
rect 13587 30209 13599 30212
rect 13541 30203 13599 30209
rect 11609 30175 11667 30181
rect 11609 30172 11621 30175
rect 11480 30144 11621 30172
rect 11480 30132 11486 30144
rect 11609 30141 11621 30144
rect 11655 30141 11667 30175
rect 11609 30135 11667 30141
rect 11885 30175 11943 30181
rect 11885 30141 11897 30175
rect 11931 30172 11943 30175
rect 13814 30172 13820 30184
rect 11931 30144 13820 30172
rect 11931 30141 11943 30144
rect 11885 30135 11943 30141
rect 13814 30132 13820 30144
rect 13872 30132 13878 30184
rect 13722 30104 13728 30116
rect 13683 30076 13728 30104
rect 13722 30064 13728 30076
rect 13780 30064 13786 30116
rect 13924 30104 13952 30212
rect 14458 30200 14464 30212
rect 14516 30200 14522 30252
rect 14737 30243 14795 30249
rect 14737 30209 14749 30243
rect 14783 30240 14795 30243
rect 15197 30243 15255 30249
rect 15197 30240 15209 30243
rect 14783 30212 15209 30240
rect 14783 30209 14795 30212
rect 14737 30203 14795 30209
rect 15197 30209 15209 30212
rect 15243 30209 15255 30243
rect 15197 30203 15255 30209
rect 15473 30243 15531 30249
rect 15473 30209 15485 30243
rect 15519 30240 15531 30243
rect 16574 30240 16580 30252
rect 15519 30212 16580 30240
rect 15519 30209 15531 30212
rect 15473 30203 15531 30209
rect 13998 30132 14004 30184
rect 14056 30172 14062 30184
rect 14752 30172 14780 30203
rect 14056 30144 14780 30172
rect 14056 30132 14062 30144
rect 15289 30107 15347 30113
rect 15289 30104 15301 30107
rect 13924 30076 15301 30104
rect 15289 30073 15301 30076
rect 15335 30073 15347 30107
rect 15289 30067 15347 30073
rect 1394 29996 1400 30048
rect 1452 30036 1458 30048
rect 1765 30039 1823 30045
rect 1765 30036 1777 30039
rect 1452 30008 1777 30036
rect 1452 29996 1458 30008
rect 1765 30005 1777 30008
rect 1811 30005 1823 30039
rect 2314 30036 2320 30048
rect 2275 30008 2320 30036
rect 1765 29999 1823 30005
rect 2314 29996 2320 30008
rect 2372 29996 2378 30048
rect 9125 30039 9183 30045
rect 9125 30005 9137 30039
rect 9171 30036 9183 30039
rect 9306 30036 9312 30048
rect 9171 30008 9312 30036
rect 9171 30005 9183 30008
rect 9125 29999 9183 30005
rect 9306 29996 9312 30008
rect 9364 29996 9370 30048
rect 13078 30036 13084 30048
rect 13039 30008 13084 30036
rect 13078 29996 13084 30008
rect 13136 29996 13142 30048
rect 14458 29996 14464 30048
rect 14516 30036 14522 30048
rect 15488 30036 15516 30203
rect 16574 30200 16580 30212
rect 16632 30200 16638 30252
rect 16853 30243 16911 30249
rect 16853 30209 16865 30243
rect 16899 30209 16911 30243
rect 16853 30203 16911 30209
rect 16868 30172 16896 30203
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 17494 30240 17500 30252
rect 17000 30212 17045 30240
rect 17455 30212 17500 30240
rect 17000 30200 17006 30212
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 18141 30243 18199 30249
rect 18141 30209 18153 30243
rect 18187 30240 18199 30243
rect 19426 30240 19432 30252
rect 18187 30212 19432 30240
rect 18187 30209 18199 30212
rect 18141 30203 18199 30209
rect 19426 30200 19432 30212
rect 19484 30200 19490 30252
rect 20990 30200 20996 30252
rect 21048 30240 21054 30252
rect 22940 30249 22968 30280
rect 26326 30268 26332 30280
rect 26384 30268 26390 30320
rect 31312 30255 31340 30348
rect 31386 30336 31392 30388
rect 31444 30376 31450 30388
rect 31444 30348 31524 30376
rect 31444 30336 31450 30348
rect 21085 30243 21143 30249
rect 21085 30240 21097 30243
rect 21048 30212 21097 30240
rect 21048 30200 21054 30212
rect 21085 30209 21097 30212
rect 21131 30209 21143 30243
rect 21085 30203 21143 30209
rect 22925 30243 22983 30249
rect 22925 30209 22937 30243
rect 22971 30209 22983 30243
rect 22925 30203 22983 30209
rect 23014 30200 23020 30252
rect 23072 30240 23078 30252
rect 23181 30243 23239 30249
rect 23181 30240 23193 30243
rect 23072 30212 23193 30240
rect 23072 30200 23078 30212
rect 23181 30209 23193 30212
rect 23227 30209 23239 30243
rect 23181 30203 23239 30209
rect 23566 30200 23572 30252
rect 23624 30240 23630 30252
rect 24857 30243 24915 30249
rect 23624 30212 23980 30240
rect 23624 30200 23630 30212
rect 17402 30172 17408 30184
rect 16592 30144 17408 30172
rect 16592 30116 16620 30144
rect 17402 30132 17408 30144
rect 17460 30132 17466 30184
rect 18414 30172 18420 30184
rect 18375 30144 18420 30172
rect 18414 30132 18420 30144
rect 18472 30132 18478 30184
rect 23952 30172 23980 30212
rect 24857 30209 24869 30243
rect 24903 30240 24915 30243
rect 25038 30240 25044 30252
rect 24903 30212 25044 30240
rect 24903 30209 24915 30212
rect 24857 30203 24915 30209
rect 25038 30200 25044 30212
rect 25096 30200 25102 30252
rect 25406 30200 25412 30252
rect 25464 30240 25470 30252
rect 25501 30243 25559 30249
rect 25501 30240 25513 30243
rect 25464 30212 25513 30240
rect 25464 30200 25470 30212
rect 25501 30209 25513 30212
rect 25547 30209 25559 30243
rect 25501 30203 25559 30209
rect 25685 30243 25743 30249
rect 25685 30209 25697 30243
rect 25731 30209 25743 30243
rect 25685 30203 25743 30209
rect 25700 30172 25728 30203
rect 30926 30200 30932 30252
rect 30984 30240 30990 30252
rect 31294 30249 31352 30255
rect 31185 30243 31243 30249
rect 31185 30240 31197 30243
rect 30984 30212 31197 30240
rect 30984 30200 30990 30212
rect 31185 30209 31197 30212
rect 31231 30209 31243 30243
rect 31294 30215 31306 30249
rect 31340 30215 31352 30249
rect 31294 30209 31352 30215
rect 31410 30243 31468 30249
rect 31410 30209 31422 30243
rect 31456 30240 31468 30243
rect 31496 30240 31524 30348
rect 33594 30308 33600 30320
rect 33555 30280 33600 30308
rect 33594 30268 33600 30280
rect 33652 30268 33658 30320
rect 31456 30212 31524 30240
rect 31573 30243 31631 30249
rect 31456 30209 31468 30212
rect 31185 30203 31243 30209
rect 31410 30203 31468 30209
rect 31573 30209 31585 30243
rect 31619 30209 31631 30243
rect 31573 30203 31631 30209
rect 23952 30144 25728 30172
rect 25774 30132 25780 30184
rect 25832 30172 25838 30184
rect 29270 30172 29276 30184
rect 25832 30144 29276 30172
rect 25832 30132 25838 30144
rect 29270 30132 29276 30144
rect 29328 30132 29334 30184
rect 31588 30172 31616 30203
rect 31662 30200 31668 30252
rect 31720 30240 31726 30252
rect 31938 30240 31944 30252
rect 31720 30212 31944 30240
rect 31720 30200 31726 30212
rect 31938 30200 31944 30212
rect 31996 30200 32002 30252
rect 32122 30240 32128 30252
rect 32083 30212 32128 30240
rect 32122 30200 32128 30212
rect 32180 30200 32186 30252
rect 32306 30240 32312 30252
rect 32267 30212 32312 30240
rect 32306 30200 32312 30212
rect 32364 30200 32370 30252
rect 33226 30200 33232 30252
rect 33284 30240 33290 30252
rect 33413 30243 33471 30249
rect 33413 30240 33425 30243
rect 33284 30212 33425 30240
rect 33284 30200 33290 30212
rect 33413 30209 33425 30212
rect 33459 30209 33471 30243
rect 33413 30203 33471 30209
rect 32493 30175 32551 30181
rect 32493 30172 32505 30175
rect 31588 30144 32505 30172
rect 32493 30141 32505 30144
rect 32539 30141 32551 30175
rect 32493 30135 32551 30141
rect 35253 30175 35311 30181
rect 35253 30141 35265 30175
rect 35299 30172 35311 30175
rect 35434 30172 35440 30184
rect 35299 30144 35440 30172
rect 35299 30141 35311 30144
rect 35253 30135 35311 30141
rect 35434 30132 35440 30144
rect 35492 30132 35498 30184
rect 16574 30064 16580 30116
rect 16632 30064 16638 30116
rect 16669 30107 16727 30113
rect 16669 30073 16681 30107
rect 16715 30104 16727 30107
rect 16758 30104 16764 30116
rect 16715 30076 16764 30104
rect 16715 30073 16727 30076
rect 16669 30067 16727 30073
rect 16758 30064 16764 30076
rect 16816 30064 16822 30116
rect 35526 30104 35532 30116
rect 25792 30076 35532 30104
rect 14516 30008 15516 30036
rect 17589 30039 17647 30045
rect 14516 29996 14522 30008
rect 17589 30005 17601 30039
rect 17635 30036 17647 30039
rect 18046 30036 18052 30048
rect 17635 30008 18052 30036
rect 17635 30005 17647 30008
rect 17589 29999 17647 30005
rect 18046 29996 18052 30008
rect 18104 29996 18110 30048
rect 18138 29996 18144 30048
rect 18196 30036 18202 30048
rect 19521 30039 19579 30045
rect 19521 30036 19533 30039
rect 18196 30008 19533 30036
rect 18196 29996 18202 30008
rect 19521 30005 19533 30008
rect 19567 30036 19579 30039
rect 22738 30036 22744 30048
rect 19567 30008 22744 30036
rect 19567 30005 19579 30008
rect 19521 29999 19579 30005
rect 22738 29996 22744 30008
rect 22796 29996 22802 30048
rect 24302 30036 24308 30048
rect 24263 30008 24308 30036
rect 24302 29996 24308 30008
rect 24360 29996 24366 30048
rect 25038 29996 25044 30048
rect 25096 30036 25102 30048
rect 25792 30036 25820 30076
rect 35526 30064 35532 30076
rect 35584 30064 35590 30116
rect 25096 30008 25820 30036
rect 30929 30039 30987 30045
rect 25096 29996 25102 30008
rect 30929 30005 30941 30039
rect 30975 30036 30987 30039
rect 31846 30036 31852 30048
rect 30975 30008 31852 30036
rect 30975 30005 30987 30008
rect 30929 29999 30987 30005
rect 31846 29996 31852 30008
rect 31904 29996 31910 30048
rect 31938 29996 31944 30048
rect 31996 30036 32002 30048
rect 32306 30036 32312 30048
rect 31996 30008 32312 30036
rect 31996 29996 32002 30008
rect 32306 29996 32312 30008
rect 32364 29996 32370 30048
rect 1104 29946 48852 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 48852 29946
rect 1104 29872 48852 29894
rect 10318 29832 10324 29844
rect 10279 29804 10324 29832
rect 10318 29792 10324 29804
rect 10376 29792 10382 29844
rect 10962 29792 10968 29844
rect 11020 29832 11026 29844
rect 14093 29835 14151 29841
rect 14093 29832 14105 29835
rect 11020 29804 14105 29832
rect 11020 29792 11026 29804
rect 14093 29801 14105 29804
rect 14139 29801 14151 29835
rect 18138 29832 18144 29844
rect 14093 29795 14151 29801
rect 14476 29804 18144 29832
rect 6362 29724 6368 29776
rect 6420 29764 6426 29776
rect 14476 29764 14504 29804
rect 6420 29736 14504 29764
rect 14553 29767 14611 29773
rect 6420 29724 6426 29736
rect 14553 29733 14565 29767
rect 14599 29733 14611 29767
rect 14553 29727 14611 29733
rect 1394 29696 1400 29708
rect 1355 29668 1400 29696
rect 1394 29656 1400 29668
rect 1452 29656 1458 29708
rect 1581 29699 1639 29705
rect 1581 29665 1593 29699
rect 1627 29696 1639 29699
rect 2314 29696 2320 29708
rect 1627 29668 2320 29696
rect 1627 29665 1639 29668
rect 1581 29659 1639 29665
rect 2314 29656 2320 29668
rect 2372 29656 2378 29708
rect 2774 29656 2780 29708
rect 2832 29696 2838 29708
rect 10965 29699 11023 29705
rect 2832 29668 2877 29696
rect 2832 29656 2838 29668
rect 10965 29665 10977 29699
rect 11011 29696 11023 29699
rect 11790 29696 11796 29708
rect 11011 29668 11192 29696
rect 11703 29668 11796 29696
rect 11011 29665 11023 29668
rect 10965 29659 11023 29665
rect 9493 29631 9551 29637
rect 9493 29597 9505 29631
rect 9539 29628 9551 29631
rect 10042 29628 10048 29640
rect 9539 29600 10048 29628
rect 9539 29597 9551 29600
rect 9493 29591 9551 29597
rect 10042 29588 10048 29600
rect 10100 29588 10106 29640
rect 10594 29628 10600 29640
rect 10555 29600 10600 29628
rect 10594 29588 10600 29600
rect 10652 29588 10658 29640
rect 11057 29631 11115 29637
rect 11057 29597 11069 29631
rect 11103 29597 11115 29631
rect 11164 29628 11192 29668
rect 11790 29656 11796 29668
rect 11848 29696 11854 29708
rect 13722 29696 13728 29708
rect 11848 29668 13728 29696
rect 11848 29656 11854 29668
rect 13722 29656 13728 29668
rect 13780 29656 13786 29708
rect 13906 29656 13912 29708
rect 13964 29696 13970 29708
rect 14185 29699 14243 29705
rect 14185 29696 14197 29699
rect 13964 29668 14197 29696
rect 13964 29656 13970 29668
rect 14185 29665 14197 29668
rect 14231 29665 14243 29699
rect 14185 29659 14243 29665
rect 11330 29628 11336 29640
rect 11164 29600 11336 29628
rect 11057 29591 11115 29597
rect 9674 29560 9680 29572
rect 9635 29532 9680 29560
rect 9674 29520 9680 29532
rect 9732 29520 9738 29572
rect 9861 29563 9919 29569
rect 9861 29529 9873 29563
rect 9907 29560 9919 29563
rect 10689 29563 10747 29569
rect 10689 29560 10701 29563
rect 9907 29532 10701 29560
rect 9907 29529 9919 29532
rect 9861 29523 9919 29529
rect 10689 29529 10701 29532
rect 10735 29529 10747 29563
rect 11072 29560 11100 29591
rect 11330 29588 11336 29600
rect 11388 29628 11394 29640
rect 11517 29631 11575 29637
rect 11517 29628 11529 29631
rect 11388 29600 11529 29628
rect 11388 29588 11394 29600
rect 11517 29597 11529 29600
rect 11563 29597 11575 29631
rect 14369 29631 14427 29637
rect 14369 29628 14381 29631
rect 11517 29591 11575 29597
rect 12406 29600 14381 29628
rect 11422 29560 11428 29572
rect 11072 29532 11428 29560
rect 10689 29523 10747 29529
rect 11422 29520 11428 29532
rect 11480 29520 11486 29572
rect 10134 29452 10140 29504
rect 10192 29492 10198 29504
rect 10781 29495 10839 29501
rect 10781 29492 10793 29495
rect 10192 29464 10793 29492
rect 10192 29452 10198 29464
rect 10781 29461 10793 29464
rect 10827 29461 10839 29495
rect 10781 29455 10839 29461
rect 10870 29452 10876 29504
rect 10928 29492 10934 29504
rect 12406 29492 12434 29600
rect 14369 29597 14381 29600
rect 14415 29597 14427 29631
rect 14568 29628 14596 29727
rect 17678 29724 17684 29776
rect 17736 29724 17742 29776
rect 15197 29631 15255 29637
rect 15197 29628 15209 29631
rect 14568 29600 15209 29628
rect 14369 29591 14427 29597
rect 15197 29597 15209 29600
rect 15243 29597 15255 29631
rect 15197 29591 15255 29597
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29628 15439 29631
rect 17402 29628 17408 29640
rect 15427 29600 17408 29628
rect 15427 29597 15439 29600
rect 15381 29591 15439 29597
rect 17402 29588 17408 29600
rect 17460 29588 17466 29640
rect 17696 29637 17724 29724
rect 17788 29705 17816 29804
rect 18138 29792 18144 29804
rect 18196 29792 18202 29844
rect 18233 29835 18291 29841
rect 18233 29801 18245 29835
rect 18279 29832 18291 29835
rect 18414 29832 18420 29844
rect 18279 29804 18420 29832
rect 18279 29801 18291 29804
rect 18233 29795 18291 29801
rect 18414 29792 18420 29804
rect 18472 29792 18478 29844
rect 18506 29792 18512 29844
rect 18564 29832 18570 29844
rect 23750 29832 23756 29844
rect 18564 29804 23756 29832
rect 18564 29792 18570 29804
rect 23750 29792 23756 29804
rect 23808 29792 23814 29844
rect 25406 29792 25412 29844
rect 25464 29832 25470 29844
rect 27617 29835 27675 29841
rect 27617 29832 27629 29835
rect 25464 29804 27629 29832
rect 25464 29792 25470 29804
rect 27617 29801 27629 29804
rect 27663 29801 27675 29835
rect 27617 29795 27675 29801
rect 32122 29792 32128 29844
rect 32180 29832 32186 29844
rect 33137 29835 33195 29841
rect 33137 29832 33149 29835
rect 32180 29804 33149 29832
rect 32180 29792 32186 29804
rect 33137 29801 33149 29804
rect 33183 29832 33195 29835
rect 34514 29832 34520 29844
rect 33183 29804 34520 29832
rect 33183 29801 33195 29804
rect 33137 29795 33195 29801
rect 34514 29792 34520 29804
rect 34572 29792 34578 29844
rect 22738 29724 22744 29776
rect 22796 29764 22802 29776
rect 25774 29764 25780 29776
rect 22796 29736 25780 29764
rect 22796 29724 22802 29736
rect 25774 29724 25780 29736
rect 25832 29724 25838 29776
rect 31662 29764 31668 29776
rect 28184 29736 31668 29764
rect 28184 29708 28212 29736
rect 31662 29724 31668 29736
rect 31720 29724 31726 29776
rect 17773 29699 17831 29705
rect 17773 29665 17785 29699
rect 17819 29665 17831 29699
rect 17773 29659 17831 29665
rect 17865 29699 17923 29705
rect 17865 29665 17877 29699
rect 17911 29696 17923 29699
rect 19242 29696 19248 29708
rect 17911 29668 19248 29696
rect 17911 29665 17923 29668
rect 17865 29659 17923 29665
rect 19242 29656 19248 29668
rect 19300 29656 19306 29708
rect 27338 29656 27344 29708
rect 27396 29696 27402 29708
rect 28077 29699 28135 29705
rect 28077 29696 28089 29699
rect 27396 29668 28089 29696
rect 27396 29656 27402 29668
rect 28077 29665 28089 29668
rect 28123 29665 28135 29699
rect 28077 29659 28135 29665
rect 28166 29656 28172 29708
rect 28224 29696 28230 29708
rect 28224 29668 28269 29696
rect 28224 29656 28230 29668
rect 28442 29656 28448 29708
rect 28500 29696 28506 29708
rect 28500 29668 31156 29696
rect 28500 29656 28506 29668
rect 17497 29631 17555 29637
rect 17497 29597 17509 29631
rect 17543 29628 17555 29631
rect 17685 29631 17743 29637
rect 17543 29600 17623 29628
rect 17543 29597 17555 29600
rect 17497 29591 17555 29597
rect 14093 29563 14151 29569
rect 14093 29529 14105 29563
rect 14139 29560 14151 29563
rect 14274 29560 14280 29572
rect 14139 29532 14280 29560
rect 14139 29529 14151 29532
rect 14093 29523 14151 29529
rect 14274 29520 14280 29532
rect 14332 29520 14338 29572
rect 15838 29560 15844 29572
rect 15799 29532 15844 29560
rect 15838 29520 15844 29532
rect 15896 29520 15902 29572
rect 16022 29560 16028 29572
rect 15983 29532 16028 29560
rect 16022 29520 16028 29532
rect 16080 29520 16086 29572
rect 15286 29492 15292 29504
rect 10928 29464 12434 29492
rect 15247 29464 15292 29492
rect 10928 29452 10934 29464
rect 15286 29452 15292 29464
rect 15344 29452 15350 29504
rect 15930 29452 15936 29504
rect 15988 29492 15994 29504
rect 16209 29495 16267 29501
rect 16209 29492 16221 29495
rect 15988 29464 16221 29492
rect 15988 29452 15994 29464
rect 16209 29461 16221 29464
rect 16255 29461 16267 29495
rect 16209 29455 16267 29461
rect 16298 29452 16304 29504
rect 16356 29492 16362 29504
rect 17595 29492 17623 29600
rect 17685 29597 17697 29631
rect 17731 29597 17743 29631
rect 18046 29628 18052 29640
rect 18007 29600 18052 29628
rect 17685 29591 17743 29597
rect 18046 29588 18052 29600
rect 18104 29588 18110 29640
rect 19426 29588 19432 29640
rect 19484 29628 19490 29640
rect 20717 29631 20775 29637
rect 20717 29628 20729 29631
rect 19484 29600 20729 29628
rect 19484 29588 19490 29600
rect 20717 29597 20729 29600
rect 20763 29597 20775 29631
rect 20717 29591 20775 29597
rect 20806 29588 20812 29640
rect 20864 29628 20870 29640
rect 20973 29631 21031 29637
rect 20973 29628 20985 29631
rect 20864 29600 20985 29628
rect 20864 29588 20870 29600
rect 20973 29597 20985 29600
rect 21019 29597 21031 29631
rect 20973 29591 21031 29597
rect 25777 29631 25835 29637
rect 25777 29597 25789 29631
rect 25823 29628 25835 29631
rect 26326 29628 26332 29640
rect 25823 29600 26332 29628
rect 25823 29597 25835 29600
rect 25777 29591 25835 29597
rect 26326 29588 26332 29600
rect 26384 29588 26390 29640
rect 27246 29588 27252 29640
rect 27304 29628 27310 29640
rect 27798 29628 27804 29640
rect 27304 29600 27804 29628
rect 27304 29588 27310 29600
rect 27798 29588 27804 29600
rect 27856 29628 27862 29640
rect 30926 29628 30932 29640
rect 27856 29600 30932 29628
rect 27856 29588 27862 29600
rect 30926 29588 30932 29600
rect 30984 29588 30990 29640
rect 31128 29637 31156 29668
rect 31202 29656 31208 29708
rect 31260 29696 31266 29708
rect 31754 29696 31760 29708
rect 31260 29668 31760 29696
rect 31260 29656 31266 29668
rect 31754 29656 31760 29668
rect 31812 29696 31818 29708
rect 35526 29696 35532 29708
rect 31812 29668 31905 29696
rect 35487 29668 35532 29696
rect 31812 29656 31818 29668
rect 35526 29656 35532 29668
rect 35584 29656 35590 29708
rect 42794 29656 42800 29708
rect 42852 29696 42858 29708
rect 47581 29699 47639 29705
rect 47581 29696 47593 29699
rect 42852 29668 47593 29696
rect 42852 29656 42858 29668
rect 47581 29665 47593 29668
rect 47627 29665 47639 29699
rect 47581 29659 47639 29665
rect 31021 29631 31079 29637
rect 31021 29597 31033 29631
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 31113 29631 31171 29637
rect 31113 29597 31125 29631
rect 31159 29597 31171 29631
rect 31113 29591 31171 29597
rect 31297 29631 31355 29637
rect 31297 29597 31309 29631
rect 31343 29628 31355 29631
rect 31343 29600 31754 29628
rect 31343 29597 31355 29600
rect 31297 29591 31355 29597
rect 19334 29520 19340 29572
rect 19392 29560 19398 29572
rect 19705 29563 19763 29569
rect 19705 29560 19717 29563
rect 19392 29532 19717 29560
rect 19392 29520 19398 29532
rect 19705 29529 19717 29532
rect 19751 29560 19763 29563
rect 20622 29560 20628 29572
rect 19751 29532 20628 29560
rect 19751 29529 19763 29532
rect 19705 29523 19763 29529
rect 20622 29520 20628 29532
rect 20680 29520 20686 29572
rect 25590 29520 25596 29572
rect 25648 29560 25654 29572
rect 26022 29563 26080 29569
rect 26022 29560 26034 29563
rect 25648 29532 26034 29560
rect 25648 29520 25654 29532
rect 26022 29529 26034 29532
rect 26068 29529 26080 29563
rect 31036 29560 31064 29591
rect 26022 29523 26080 29529
rect 26160 29532 31064 29560
rect 31128 29560 31156 29591
rect 31386 29560 31392 29572
rect 31128 29532 31392 29560
rect 18690 29492 18696 29504
rect 16356 29464 18696 29492
rect 16356 29452 16362 29464
rect 18690 29452 18696 29464
rect 18748 29492 18754 29504
rect 19797 29495 19855 29501
rect 19797 29492 19809 29495
rect 18748 29464 19809 29492
rect 18748 29452 18754 29464
rect 19797 29461 19809 29464
rect 19843 29461 19855 29495
rect 19797 29455 19855 29461
rect 22097 29495 22155 29501
rect 22097 29461 22109 29495
rect 22143 29492 22155 29495
rect 22186 29492 22192 29504
rect 22143 29464 22192 29492
rect 22143 29461 22155 29464
rect 22097 29455 22155 29461
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 24302 29452 24308 29504
rect 24360 29492 24366 29504
rect 26160 29492 26188 29532
rect 31386 29520 31392 29532
rect 31444 29520 31450 29572
rect 31726 29560 31754 29600
rect 31846 29588 31852 29640
rect 31904 29628 31910 29640
rect 32013 29631 32071 29637
rect 32013 29628 32025 29631
rect 31904 29600 32025 29628
rect 31904 29588 31910 29600
rect 32013 29597 32025 29600
rect 32059 29597 32071 29631
rect 32013 29591 32071 29597
rect 33502 29588 33508 29640
rect 33560 29628 33566 29640
rect 33597 29631 33655 29637
rect 33597 29628 33609 29631
rect 33560 29600 33609 29628
rect 33560 29588 33566 29600
rect 33597 29597 33609 29600
rect 33643 29597 33655 29631
rect 33597 29591 33655 29597
rect 33962 29588 33968 29640
rect 34020 29628 34026 29640
rect 34606 29628 34612 29640
rect 34020 29600 34612 29628
rect 34020 29588 34026 29600
rect 34606 29588 34612 29600
rect 34664 29628 34670 29640
rect 34701 29631 34759 29637
rect 34701 29628 34713 29631
rect 34664 29600 34713 29628
rect 34664 29588 34670 29600
rect 34701 29597 34713 29600
rect 34747 29597 34759 29631
rect 47302 29628 47308 29640
rect 47263 29600 47308 29628
rect 34701 29591 34759 29597
rect 47302 29588 47308 29600
rect 47360 29588 47366 29640
rect 32214 29560 32220 29572
rect 31726 29532 32220 29560
rect 32214 29520 32220 29532
rect 32272 29520 32278 29572
rect 35710 29560 35716 29572
rect 35671 29532 35716 29560
rect 35710 29520 35716 29532
rect 35768 29520 35774 29572
rect 37369 29563 37427 29569
rect 37369 29529 37381 29563
rect 37415 29560 37427 29563
rect 46842 29560 46848 29572
rect 37415 29532 46848 29560
rect 37415 29529 37427 29532
rect 37369 29523 37427 29529
rect 46842 29520 46848 29532
rect 46900 29520 46906 29572
rect 24360 29464 26188 29492
rect 27157 29495 27215 29501
rect 24360 29452 24366 29464
rect 27157 29461 27169 29495
rect 27203 29492 27215 29495
rect 27706 29492 27712 29504
rect 27203 29464 27712 29492
rect 27203 29461 27215 29464
rect 27157 29455 27215 29461
rect 27706 29452 27712 29464
rect 27764 29492 27770 29504
rect 27985 29495 28043 29501
rect 27985 29492 27997 29495
rect 27764 29464 27997 29492
rect 27764 29452 27770 29464
rect 27985 29461 27997 29464
rect 28031 29461 28043 29495
rect 27985 29455 28043 29461
rect 30653 29495 30711 29501
rect 30653 29461 30665 29495
rect 30699 29492 30711 29495
rect 32122 29492 32128 29504
rect 30699 29464 32128 29492
rect 30699 29461 30711 29464
rect 30653 29455 30711 29461
rect 32122 29452 32128 29464
rect 32180 29452 32186 29504
rect 33686 29492 33692 29504
rect 33647 29464 33692 29492
rect 33686 29452 33692 29464
rect 33744 29452 33750 29504
rect 34790 29492 34796 29504
rect 34751 29464 34796 29492
rect 34790 29452 34796 29464
rect 34848 29452 34854 29504
rect 1104 29402 48852 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 48852 29402
rect 1104 29328 48852 29350
rect 9950 29288 9956 29300
rect 9911 29260 9956 29288
rect 9950 29248 9956 29260
rect 10008 29248 10014 29300
rect 10042 29248 10048 29300
rect 10100 29288 10106 29300
rect 10873 29291 10931 29297
rect 10873 29288 10885 29291
rect 10100 29260 10885 29288
rect 10100 29248 10106 29260
rect 10873 29257 10885 29260
rect 10919 29257 10931 29291
rect 10873 29251 10931 29257
rect 11701 29291 11759 29297
rect 11701 29257 11713 29291
rect 11747 29288 11759 29291
rect 11790 29288 11796 29300
rect 11747 29260 11796 29288
rect 11747 29257 11759 29260
rect 11701 29251 11759 29257
rect 11790 29248 11796 29260
rect 11848 29248 11854 29300
rect 14458 29248 14464 29300
rect 14516 29288 14522 29300
rect 14737 29291 14795 29297
rect 14737 29288 14749 29291
rect 14516 29260 14749 29288
rect 14516 29248 14522 29260
rect 14737 29257 14749 29260
rect 14783 29257 14795 29291
rect 14737 29251 14795 29257
rect 15286 29248 15292 29300
rect 15344 29288 15350 29300
rect 15344 29260 22094 29288
rect 15344 29248 15350 29260
rect 9214 29180 9220 29232
rect 9272 29220 9278 29232
rect 10505 29223 10563 29229
rect 10505 29220 10517 29223
rect 9272 29192 10517 29220
rect 9272 29180 9278 29192
rect 10505 29189 10517 29192
rect 10551 29189 10563 29223
rect 10505 29183 10563 29189
rect 10721 29223 10779 29229
rect 10721 29189 10733 29223
rect 10767 29220 10779 29223
rect 12980 29223 13038 29229
rect 10767 29192 11836 29220
rect 10767 29189 10779 29192
rect 10721 29183 10779 29189
rect 2317 29155 2375 29161
rect 2317 29121 2329 29155
rect 2363 29152 2375 29155
rect 2682 29152 2688 29164
rect 2363 29124 2688 29152
rect 2363 29121 2375 29124
rect 2317 29115 2375 29121
rect 2682 29112 2688 29124
rect 2740 29112 2746 29164
rect 2958 29152 2964 29164
rect 2919 29124 2964 29152
rect 2958 29112 2964 29124
rect 3016 29112 3022 29164
rect 9861 29155 9919 29161
rect 9861 29121 9873 29155
rect 9907 29121 9919 29155
rect 10042 29152 10048 29164
rect 10003 29124 10048 29152
rect 9861 29115 9919 29121
rect 9876 29084 9904 29115
rect 10042 29112 10048 29124
rect 10100 29112 10106 29164
rect 10520 29152 10548 29183
rect 11808 29161 11836 29192
rect 12980 29189 12992 29223
rect 13026 29220 13038 29223
rect 13078 29220 13084 29232
rect 13026 29192 13084 29220
rect 13026 29189 13038 29192
rect 12980 29183 13038 29189
rect 13078 29180 13084 29192
rect 13136 29180 13142 29232
rect 16482 29220 16488 29232
rect 14568 29192 16488 29220
rect 11517 29155 11575 29161
rect 11517 29152 11529 29155
rect 10520 29124 11529 29152
rect 11517 29121 11529 29124
rect 11563 29152 11575 29155
rect 11793 29155 11851 29161
rect 11563 29124 11652 29152
rect 11563 29121 11575 29124
rect 11517 29115 11575 29121
rect 9876 29056 11560 29084
rect 11532 29025 11560 29056
rect 11517 29019 11575 29025
rect 11517 28985 11529 29019
rect 11563 28985 11575 29019
rect 11624 29016 11652 29124
rect 11793 29121 11805 29155
rect 11839 29152 11851 29155
rect 12710 29152 12716 29164
rect 11839 29124 12572 29152
rect 12671 29124 12716 29152
rect 11839 29121 11851 29124
rect 11793 29115 11851 29121
rect 12544 29084 12572 29124
rect 12710 29112 12716 29124
rect 12768 29112 12774 29164
rect 14568 29152 14596 29192
rect 15764 29161 15792 29192
rect 16482 29180 16488 29192
rect 16540 29180 16546 29232
rect 19426 29220 19432 29232
rect 16684 29192 19432 29220
rect 12820 29124 14596 29152
rect 14645 29155 14703 29161
rect 12618 29084 12624 29096
rect 12544 29056 12624 29084
rect 12618 29044 12624 29056
rect 12676 29044 12682 29096
rect 12820 29084 12848 29124
rect 14645 29121 14657 29155
rect 14691 29121 14703 29155
rect 14645 29115 14703 29121
rect 15749 29155 15807 29161
rect 15749 29121 15761 29155
rect 15795 29121 15807 29155
rect 15749 29115 15807 29121
rect 15841 29155 15899 29161
rect 15841 29121 15853 29155
rect 15887 29121 15899 29155
rect 15841 29115 15899 29121
rect 12728 29056 12848 29084
rect 12728 29016 12756 29056
rect 14090 29016 14096 29028
rect 11624 28988 12756 29016
rect 14003 28988 14096 29016
rect 11517 28979 11575 28985
rect 14090 28976 14096 28988
rect 14148 29016 14154 29028
rect 14660 29016 14688 29115
rect 15654 29044 15660 29096
rect 15712 29084 15718 29096
rect 15856 29084 15884 29115
rect 15930 29112 15936 29164
rect 15988 29152 15994 29164
rect 15988 29124 16033 29152
rect 15988 29112 15994 29124
rect 16114 29112 16120 29164
rect 16172 29152 16178 29164
rect 16298 29152 16304 29164
rect 16172 29124 16304 29152
rect 16172 29112 16178 29124
rect 16298 29112 16304 29124
rect 16356 29112 16362 29164
rect 16684 29161 16712 29192
rect 19426 29180 19432 29192
rect 19484 29180 19490 29232
rect 16669 29155 16727 29161
rect 16669 29121 16681 29155
rect 16715 29121 16727 29155
rect 16925 29155 16983 29161
rect 16925 29152 16937 29155
rect 16669 29115 16727 29121
rect 16776 29124 16937 29152
rect 16776 29084 16804 29124
rect 16925 29121 16937 29124
rect 16971 29121 16983 29155
rect 16925 29115 16983 29121
rect 17310 29112 17316 29164
rect 17368 29152 17374 29164
rect 17862 29152 17868 29164
rect 17368 29124 17868 29152
rect 17368 29112 17374 29124
rect 17862 29112 17868 29124
rect 17920 29152 17926 29164
rect 19061 29155 19119 29161
rect 19061 29152 19073 29155
rect 17920 29124 19073 29152
rect 17920 29112 17926 29124
rect 19061 29121 19073 29124
rect 19107 29121 19119 29155
rect 19061 29115 19119 29121
rect 19245 29155 19303 29161
rect 19245 29121 19257 29155
rect 19291 29152 19303 29155
rect 21082 29152 21088 29164
rect 19291 29124 21088 29152
rect 19291 29121 19303 29124
rect 19245 29115 19303 29121
rect 21082 29112 21088 29124
rect 21140 29112 21146 29164
rect 22066 29152 22094 29260
rect 22186 29248 22192 29300
rect 22244 29288 22250 29300
rect 22244 29260 29316 29288
rect 22244 29248 22250 29260
rect 23566 29220 23572 29232
rect 23527 29192 23572 29220
rect 23566 29180 23572 29192
rect 23624 29180 23630 29232
rect 23750 29180 23756 29232
rect 23808 29220 23814 29232
rect 28442 29220 28448 29232
rect 23808 29192 28448 29220
rect 23808 29180 23814 29192
rect 28442 29180 28448 29192
rect 28500 29180 28506 29232
rect 28994 29220 29000 29232
rect 28644 29192 29000 29220
rect 28644 29161 28672 29192
rect 28994 29180 29000 29192
rect 29052 29180 29058 29232
rect 23385 29155 23443 29161
rect 23385 29152 23397 29155
rect 22066 29124 23397 29152
rect 23385 29121 23397 29124
rect 23431 29121 23443 29155
rect 25685 29155 25743 29161
rect 25685 29152 25697 29155
rect 23385 29115 23443 29121
rect 24780 29124 25697 29152
rect 15712 29056 15884 29084
rect 15948 29056 16804 29084
rect 15712 29044 15718 29056
rect 14148 28988 14688 29016
rect 14148 28976 14154 28988
rect 1854 28948 1860 28960
rect 1815 28920 1860 28948
rect 1854 28908 1860 28920
rect 1912 28908 1918 28960
rect 2406 28948 2412 28960
rect 2367 28920 2412 28948
rect 2406 28908 2412 28920
rect 2464 28908 2470 28960
rect 2866 28908 2872 28960
rect 2924 28948 2930 28960
rect 3053 28951 3111 28957
rect 3053 28948 3065 28951
rect 2924 28920 3065 28948
rect 2924 28908 2930 28920
rect 3053 28917 3065 28920
rect 3099 28917 3111 28951
rect 3053 28911 3111 28917
rect 10689 28951 10747 28957
rect 10689 28917 10701 28951
rect 10735 28948 10747 28951
rect 11238 28948 11244 28960
rect 10735 28920 11244 28948
rect 10735 28917 10747 28920
rect 10689 28911 10747 28917
rect 11238 28908 11244 28920
rect 11296 28908 11302 28960
rect 15473 28951 15531 28957
rect 15473 28917 15485 28951
rect 15519 28948 15531 28951
rect 15948 28948 15976 29056
rect 23106 29044 23112 29096
rect 23164 29084 23170 29096
rect 24780 29084 24808 29124
rect 25685 29121 25697 29124
rect 25731 29121 25743 29155
rect 25685 29115 25743 29121
rect 28629 29155 28687 29161
rect 28629 29121 28641 29155
rect 28675 29121 28687 29155
rect 28629 29115 28687 29121
rect 28896 29155 28954 29161
rect 28896 29121 28908 29155
rect 28942 29152 28954 29155
rect 29178 29152 29184 29164
rect 28942 29124 29184 29152
rect 28942 29121 28954 29124
rect 28896 29115 28954 29121
rect 29178 29112 29184 29124
rect 29236 29112 29242 29164
rect 29288 29152 29316 29260
rect 29638 29248 29644 29300
rect 29696 29288 29702 29300
rect 29822 29288 29828 29300
rect 29696 29260 29828 29288
rect 29696 29248 29702 29260
rect 29822 29248 29828 29260
rect 29880 29288 29886 29300
rect 30009 29291 30067 29297
rect 30009 29288 30021 29291
rect 29880 29260 30021 29288
rect 29880 29248 29886 29260
rect 30009 29257 30021 29260
rect 30055 29257 30067 29291
rect 30009 29251 30067 29257
rect 33410 29248 33416 29300
rect 33468 29288 33474 29300
rect 33597 29291 33655 29297
rect 33597 29288 33609 29291
rect 33468 29260 33609 29288
rect 33468 29248 33474 29260
rect 33597 29257 33609 29260
rect 33643 29257 33655 29291
rect 33597 29251 33655 29257
rect 35710 29248 35716 29300
rect 35768 29288 35774 29300
rect 37369 29291 37427 29297
rect 37369 29288 37381 29291
rect 35768 29260 37381 29288
rect 35768 29248 35774 29260
rect 37369 29257 37381 29260
rect 37415 29257 37427 29291
rect 37369 29251 37427 29257
rect 29362 29180 29368 29232
rect 29420 29220 29426 29232
rect 29420 29192 31248 29220
rect 29420 29180 29426 29192
rect 31220 29161 31248 29192
rect 32122 29180 32128 29232
rect 32180 29220 32186 29232
rect 32462 29223 32520 29229
rect 32462 29220 32474 29223
rect 32180 29192 32474 29220
rect 32180 29180 32186 29192
rect 32462 29189 32474 29192
rect 32508 29189 32520 29223
rect 37458 29220 37464 29232
rect 32462 29183 32520 29189
rect 32600 29192 37464 29220
rect 31113 29155 31171 29161
rect 31113 29152 31125 29155
rect 29288 29124 31125 29152
rect 31113 29121 31125 29124
rect 31159 29121 31171 29155
rect 31113 29115 31171 29121
rect 31205 29155 31263 29161
rect 31205 29121 31217 29155
rect 31251 29121 31263 29155
rect 31205 29115 31263 29121
rect 31297 29155 31355 29161
rect 31297 29121 31309 29155
rect 31343 29152 31355 29155
rect 31386 29152 31392 29164
rect 31343 29124 31392 29152
rect 31343 29121 31355 29124
rect 31297 29115 31355 29121
rect 31386 29112 31392 29124
rect 31444 29112 31450 29164
rect 31481 29155 31539 29161
rect 31481 29121 31493 29155
rect 31527 29121 31539 29155
rect 31481 29115 31539 29121
rect 23164 29056 24808 29084
rect 25225 29087 25283 29093
rect 23164 29044 23170 29056
rect 25225 29053 25237 29087
rect 25271 29053 25283 29087
rect 25774 29084 25780 29096
rect 25735 29056 25780 29084
rect 25225 29047 25283 29053
rect 18046 29016 18052 29028
rect 18007 28988 18052 29016
rect 18046 28976 18052 28988
rect 18104 29016 18110 29028
rect 25038 29016 25044 29028
rect 18104 28988 25044 29016
rect 18104 28976 18110 28988
rect 25038 28976 25044 28988
rect 25096 28976 25102 29028
rect 25240 29016 25268 29047
rect 25774 29044 25780 29056
rect 25832 29044 25838 29096
rect 31496 29084 31524 29115
rect 31754 29112 31760 29164
rect 31812 29152 31818 29164
rect 32217 29155 32275 29161
rect 32217 29152 32229 29155
rect 31812 29124 32229 29152
rect 31812 29112 31818 29124
rect 32217 29121 32229 29124
rect 32263 29121 32275 29155
rect 32600 29152 32628 29192
rect 37458 29180 37464 29192
rect 37516 29180 37522 29232
rect 34514 29152 34520 29164
rect 32217 29115 32275 29121
rect 32324 29124 32628 29152
rect 34475 29124 34520 29152
rect 32122 29084 32128 29096
rect 31496 29056 32128 29084
rect 32122 29044 32128 29056
rect 32180 29044 32186 29096
rect 32324 29084 32352 29124
rect 34514 29112 34520 29124
rect 34572 29112 34578 29164
rect 37274 29152 37280 29164
rect 37235 29124 37280 29152
rect 37274 29112 37280 29124
rect 37332 29112 37338 29164
rect 45830 29112 45836 29164
rect 45888 29152 45894 29164
rect 47210 29152 47216 29164
rect 45888 29124 47216 29152
rect 45888 29112 45894 29124
rect 47210 29112 47216 29124
rect 47268 29152 47274 29164
rect 47581 29155 47639 29161
rect 47581 29152 47593 29155
rect 47268 29124 47593 29152
rect 47268 29112 47274 29124
rect 47581 29121 47593 29124
rect 47627 29121 47639 29155
rect 47581 29115 47639 29121
rect 34698 29084 34704 29096
rect 32232 29056 32352 29084
rect 34659 29056 34704 29084
rect 32232 29016 32260 29056
rect 34698 29044 34704 29056
rect 34756 29044 34762 29096
rect 36354 29084 36360 29096
rect 36315 29056 36360 29084
rect 36354 29044 36360 29056
rect 36412 29044 36418 29096
rect 25240 28988 28672 29016
rect 15519 28920 15976 28948
rect 15519 28917 15531 28920
rect 15473 28911 15531 28917
rect 16574 28908 16580 28960
rect 16632 28948 16638 28960
rect 17310 28948 17316 28960
rect 16632 28920 17316 28948
rect 16632 28908 16638 28920
rect 17310 28908 17316 28920
rect 17368 28908 17374 28960
rect 19334 28908 19340 28960
rect 19392 28948 19398 28960
rect 19429 28951 19487 28957
rect 19429 28948 19441 28951
rect 19392 28920 19441 28948
rect 19392 28908 19398 28920
rect 19429 28917 19441 28920
rect 19475 28917 19487 28951
rect 19429 28911 19487 28917
rect 23290 28908 23296 28960
rect 23348 28948 23354 28960
rect 25866 28948 25872 28960
rect 23348 28920 25872 28948
rect 23348 28908 23354 28920
rect 25866 28908 25872 28920
rect 25924 28908 25930 28960
rect 28644 28948 28672 28988
rect 29564 28988 32260 29016
rect 29564 28948 29592 28988
rect 34882 28976 34888 29028
rect 34940 28976 34946 29028
rect 30834 28948 30840 28960
rect 28644 28920 29592 28948
rect 30795 28920 30840 28948
rect 30834 28908 30840 28920
rect 30892 28908 30898 28960
rect 34054 28908 34060 28960
rect 34112 28948 34118 28960
rect 34900 28948 34928 28976
rect 47026 28948 47032 28960
rect 34112 28920 34928 28948
rect 46987 28920 47032 28948
rect 34112 28908 34118 28920
rect 47026 28908 47032 28920
rect 47084 28908 47090 28960
rect 47670 28948 47676 28960
rect 47631 28920 47676 28948
rect 47670 28908 47676 28920
rect 47728 28908 47734 28960
rect 1104 28858 48852 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 48852 28858
rect 1104 28784 48852 28806
rect 10042 28744 10048 28756
rect 9232 28716 10048 28744
rect 1397 28611 1455 28617
rect 1397 28577 1409 28611
rect 1443 28608 1455 28611
rect 1854 28608 1860 28620
rect 1443 28580 1860 28608
rect 1443 28577 1455 28580
rect 1397 28571 1455 28577
rect 1854 28568 1860 28580
rect 1912 28568 1918 28620
rect 2774 28568 2780 28620
rect 2832 28608 2838 28620
rect 2832 28580 2877 28608
rect 2832 28568 2838 28580
rect 8389 28543 8447 28549
rect 8389 28509 8401 28543
rect 8435 28540 8447 28543
rect 9122 28540 9128 28552
rect 8435 28512 9128 28540
rect 8435 28509 8447 28512
rect 8389 28503 8447 28509
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 9232 28549 9260 28716
rect 10042 28704 10048 28716
rect 10100 28744 10106 28756
rect 10870 28744 10876 28756
rect 10100 28716 10876 28744
rect 10100 28704 10106 28716
rect 10870 28704 10876 28716
rect 10928 28704 10934 28756
rect 17310 28744 17316 28756
rect 17271 28716 17316 28744
rect 17310 28704 17316 28716
rect 17368 28704 17374 28756
rect 17402 28704 17408 28756
rect 17460 28744 17466 28756
rect 17497 28747 17555 28753
rect 17497 28744 17509 28747
rect 17460 28716 17509 28744
rect 17460 28704 17466 28716
rect 17497 28713 17509 28716
rect 17543 28713 17555 28747
rect 18230 28744 18236 28756
rect 17497 28707 17555 28713
rect 17604 28716 18236 28744
rect 9490 28676 9496 28688
rect 9324 28648 9496 28676
rect 9324 28549 9352 28648
rect 9490 28636 9496 28648
rect 9548 28676 9554 28688
rect 11146 28676 11152 28688
rect 9548 28648 11152 28676
rect 9548 28636 9554 28648
rect 11146 28636 11152 28648
rect 11204 28636 11210 28688
rect 11330 28636 11336 28688
rect 11388 28636 11394 28688
rect 11514 28636 11520 28688
rect 11572 28676 11578 28688
rect 11572 28648 12572 28676
rect 11572 28636 11578 28648
rect 11241 28611 11299 28617
rect 11241 28577 11253 28611
rect 11287 28608 11299 28611
rect 11348 28608 11376 28636
rect 12544 28617 12572 28648
rect 14734 28636 14740 28688
rect 14792 28676 14798 28688
rect 17604 28676 17632 28716
rect 18230 28704 18236 28716
rect 18288 28704 18294 28756
rect 20070 28704 20076 28756
rect 20128 28744 20134 28756
rect 20990 28744 20996 28756
rect 20128 28716 20996 28744
rect 20128 28704 20134 28716
rect 20990 28704 20996 28716
rect 21048 28704 21054 28756
rect 23750 28744 23756 28756
rect 23711 28716 23756 28744
rect 23750 28704 23756 28716
rect 23808 28704 23814 28756
rect 24581 28747 24639 28753
rect 24581 28713 24593 28747
rect 24627 28744 24639 28747
rect 24762 28744 24768 28756
rect 24627 28716 24768 28744
rect 24627 28713 24639 28716
rect 24581 28707 24639 28713
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 25498 28744 25504 28756
rect 25459 28716 25504 28744
rect 25498 28704 25504 28716
rect 25556 28704 25562 28756
rect 27062 28704 27068 28756
rect 27120 28744 27126 28756
rect 33226 28744 33232 28756
rect 27120 28716 33232 28744
rect 27120 28704 27126 28716
rect 33226 28704 33232 28716
rect 33284 28704 33290 28756
rect 34698 28704 34704 28756
rect 34756 28744 34762 28756
rect 34793 28747 34851 28753
rect 34793 28744 34805 28747
rect 34756 28716 34805 28744
rect 34756 28704 34762 28716
rect 34793 28713 34805 28716
rect 34839 28713 34851 28747
rect 34793 28707 34851 28713
rect 14792 28648 17632 28676
rect 14792 28636 14798 28648
rect 12529 28611 12587 28617
rect 11287 28580 12480 28608
rect 11287 28577 11299 28580
rect 11241 28571 11299 28577
rect 12452 28552 12480 28580
rect 12529 28577 12541 28611
rect 12575 28577 12587 28611
rect 12529 28571 12587 28577
rect 13998 28568 14004 28620
rect 14056 28608 14062 28620
rect 14274 28608 14280 28620
rect 14056 28580 14280 28608
rect 14056 28568 14062 28580
rect 14274 28568 14280 28580
rect 14332 28568 14338 28620
rect 14458 28608 14464 28620
rect 14419 28580 14464 28608
rect 14458 28568 14464 28580
rect 14516 28608 14522 28620
rect 15749 28611 15807 28617
rect 14516 28580 15516 28608
rect 14516 28568 14522 28580
rect 9217 28543 9275 28549
rect 9217 28509 9229 28543
rect 9263 28509 9275 28543
rect 9217 28503 9275 28509
rect 9309 28543 9367 28549
rect 9309 28509 9321 28543
rect 9355 28509 9367 28543
rect 9309 28503 9367 28509
rect 9398 28500 9404 28552
rect 9456 28540 9462 28552
rect 9456 28512 9501 28540
rect 9456 28500 9462 28512
rect 9582 28500 9588 28552
rect 9640 28540 9646 28552
rect 9640 28512 9685 28540
rect 9640 28500 9646 28512
rect 10594 28500 10600 28552
rect 10652 28540 10658 28552
rect 10873 28543 10931 28549
rect 10873 28540 10885 28543
rect 10652 28512 10885 28540
rect 10652 28500 10658 28512
rect 10873 28509 10885 28512
rect 10919 28540 10931 28543
rect 10919 28512 11284 28540
rect 10919 28509 10931 28512
rect 10873 28503 10931 28509
rect 1581 28475 1639 28481
rect 1581 28441 1593 28475
rect 1627 28472 1639 28475
rect 2406 28472 2412 28484
rect 1627 28444 2412 28472
rect 1627 28441 1639 28444
rect 1581 28435 1639 28441
rect 2406 28432 2412 28444
rect 2464 28432 2470 28484
rect 8018 28472 8024 28484
rect 7979 28444 8024 28472
rect 8018 28432 8024 28444
rect 8076 28432 8082 28484
rect 8205 28475 8263 28481
rect 8205 28441 8217 28475
rect 8251 28472 8263 28475
rect 8570 28472 8576 28484
rect 8251 28444 8576 28472
rect 8251 28441 8263 28444
rect 8205 28435 8263 28441
rect 8570 28432 8576 28444
rect 8628 28432 8634 28484
rect 10965 28475 11023 28481
rect 10965 28441 10977 28475
rect 11011 28472 11023 28475
rect 11146 28472 11152 28484
rect 11011 28444 11152 28472
rect 11011 28441 11023 28444
rect 10965 28435 11023 28441
rect 11146 28432 11152 28444
rect 11204 28432 11210 28484
rect 11256 28472 11284 28512
rect 11330 28500 11336 28552
rect 11388 28540 11394 28552
rect 12066 28540 12072 28552
rect 11388 28512 11433 28540
rect 12027 28512 12072 28540
rect 11388 28500 11394 28512
rect 12066 28500 12072 28512
rect 12124 28500 12130 28552
rect 12434 28540 12440 28552
rect 12395 28512 12440 28540
rect 12434 28500 12440 28512
rect 12492 28500 12498 28552
rect 12618 28500 12624 28552
rect 12676 28540 12682 28552
rect 12989 28543 13047 28549
rect 12989 28540 13001 28543
rect 12676 28512 13001 28540
rect 12676 28500 12682 28512
rect 12989 28509 13001 28512
rect 13035 28509 13047 28543
rect 12989 28503 13047 28509
rect 14366 28500 14372 28552
rect 14424 28540 14430 28552
rect 14553 28543 14611 28549
rect 14424 28512 14469 28540
rect 14424 28500 14430 28512
rect 14553 28509 14565 28543
rect 14599 28540 14611 28543
rect 14734 28540 14740 28552
rect 14599 28512 14740 28540
rect 14599 28509 14611 28512
rect 14553 28503 14611 28509
rect 14734 28500 14740 28512
rect 14792 28500 14798 28552
rect 12084 28472 12112 28500
rect 11256 28444 12112 28472
rect 12161 28475 12219 28481
rect 12161 28441 12173 28475
rect 12207 28472 12219 28475
rect 15488 28472 15516 28580
rect 15749 28577 15761 28611
rect 15795 28608 15807 28611
rect 15838 28608 15844 28620
rect 15795 28580 15844 28608
rect 15795 28577 15807 28580
rect 15749 28571 15807 28577
rect 15838 28568 15844 28580
rect 15896 28568 15902 28620
rect 16025 28611 16083 28617
rect 16025 28577 16037 28611
rect 16071 28608 16083 28611
rect 16574 28608 16580 28620
rect 16071 28580 16580 28608
rect 16071 28577 16083 28580
rect 16025 28571 16083 28577
rect 16574 28568 16580 28580
rect 16632 28568 16638 28620
rect 17236 28617 17264 28648
rect 18046 28636 18052 28688
rect 18104 28676 18110 28688
rect 24780 28676 24808 28704
rect 25866 28676 25872 28688
rect 18104 28648 18149 28676
rect 24780 28648 25872 28676
rect 18104 28636 18110 28648
rect 25866 28636 25872 28648
rect 25924 28636 25930 28688
rect 27246 28676 27252 28688
rect 26068 28648 27252 28676
rect 17221 28611 17279 28617
rect 17221 28577 17233 28611
rect 17267 28577 17279 28611
rect 17221 28571 17279 28577
rect 17586 28568 17592 28620
rect 17644 28608 17650 28620
rect 19426 28608 19432 28620
rect 17644 28580 18736 28608
rect 19387 28580 19432 28608
rect 17644 28568 17650 28580
rect 16482 28500 16488 28552
rect 16540 28540 16546 28552
rect 17313 28543 17371 28549
rect 17313 28540 17325 28543
rect 16540 28512 17325 28540
rect 16540 28500 16546 28512
rect 17313 28509 17325 28512
rect 17359 28509 17371 28543
rect 17313 28503 17371 28509
rect 18138 28500 18144 28552
rect 18196 28540 18202 28552
rect 18279 28543 18337 28549
rect 18279 28540 18291 28543
rect 18196 28512 18291 28540
rect 18196 28500 18202 28512
rect 18279 28509 18291 28512
rect 18325 28509 18337 28543
rect 18279 28503 18337 28509
rect 18417 28543 18475 28549
rect 18417 28509 18429 28543
rect 18463 28509 18475 28543
rect 18417 28503 18475 28509
rect 17037 28475 17095 28481
rect 17037 28472 17049 28475
rect 12207 28444 14136 28472
rect 15488 28444 17049 28472
rect 12207 28441 12219 28444
rect 12161 28435 12219 28441
rect 8478 28364 8484 28416
rect 8536 28404 8542 28416
rect 8941 28407 8999 28413
rect 8941 28404 8953 28407
rect 8536 28376 8953 28404
rect 8536 28364 8542 28376
rect 8941 28373 8953 28376
rect 8987 28373 8999 28407
rect 10594 28404 10600 28416
rect 10555 28376 10600 28404
rect 8941 28367 8999 28373
rect 10594 28364 10600 28376
rect 10652 28364 10658 28416
rect 11054 28404 11060 28416
rect 11015 28376 11060 28404
rect 11054 28364 11060 28376
rect 11112 28364 11118 28416
rect 11793 28407 11851 28413
rect 11793 28373 11805 28407
rect 11839 28404 11851 28407
rect 11882 28404 11888 28416
rect 11839 28376 11888 28404
rect 11839 28373 11851 28376
rect 11793 28367 11851 28373
rect 11882 28364 11888 28376
rect 11940 28364 11946 28416
rect 14108 28413 14136 28444
rect 17037 28441 17049 28444
rect 17083 28441 17095 28475
rect 17037 28435 17095 28441
rect 17218 28432 17224 28484
rect 17276 28472 17282 28484
rect 18432 28472 18460 28503
rect 18506 28500 18512 28552
rect 18564 28540 18570 28552
rect 18708 28549 18736 28580
rect 19426 28568 19432 28580
rect 19484 28568 19490 28620
rect 25590 28568 25596 28620
rect 25648 28608 25654 28620
rect 25685 28611 25743 28617
rect 25685 28608 25697 28611
rect 25648 28580 25697 28608
rect 25648 28568 25654 28580
rect 25685 28577 25697 28580
rect 25731 28577 25743 28611
rect 25685 28571 25743 28577
rect 18693 28543 18751 28549
rect 18564 28512 18609 28540
rect 18564 28500 18570 28512
rect 18693 28509 18705 28543
rect 18739 28540 18751 28543
rect 18782 28540 18788 28552
rect 18739 28512 18788 28540
rect 18739 28509 18751 28512
rect 18693 28503 18751 28509
rect 18782 28500 18788 28512
rect 18840 28500 18846 28552
rect 23382 28500 23388 28552
rect 23440 28540 23446 28552
rect 23569 28543 23627 28549
rect 23569 28540 23581 28543
rect 23440 28512 23581 28540
rect 23440 28500 23446 28512
rect 23569 28509 23581 28512
rect 23615 28509 23627 28543
rect 23569 28503 23627 28509
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 25130 28540 25136 28552
rect 24443 28512 25136 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 25130 28500 25136 28512
rect 25188 28500 25194 28552
rect 25409 28543 25467 28549
rect 25409 28509 25421 28543
rect 25455 28540 25467 28543
rect 26068 28540 26096 28648
rect 27246 28636 27252 28648
rect 27304 28636 27310 28688
rect 28994 28636 29000 28688
rect 29052 28676 29058 28688
rect 29546 28676 29552 28688
rect 29052 28648 29552 28676
rect 29052 28636 29058 28648
rect 29546 28636 29552 28648
rect 29604 28676 29610 28688
rect 29604 28648 31248 28676
rect 29604 28636 29610 28648
rect 31220 28620 31248 28648
rect 26421 28611 26479 28617
rect 26421 28577 26433 28611
rect 26467 28608 26479 28611
rect 28166 28608 28172 28620
rect 26467 28580 28172 28608
rect 26467 28577 26479 28580
rect 26421 28571 26479 28577
rect 28166 28568 28172 28580
rect 28224 28608 28230 28620
rect 29917 28611 29975 28617
rect 29917 28608 29929 28611
rect 28224 28580 29929 28608
rect 28224 28568 28230 28580
rect 29917 28577 29929 28580
rect 29963 28577 29975 28611
rect 29917 28571 29975 28577
rect 30098 28568 30104 28620
rect 30156 28608 30162 28620
rect 30193 28611 30251 28617
rect 30193 28608 30205 28611
rect 30156 28580 30205 28608
rect 30156 28568 30162 28580
rect 30193 28577 30205 28580
rect 30239 28577 30251 28611
rect 31202 28608 31208 28620
rect 31163 28580 31208 28608
rect 30193 28571 30251 28577
rect 31202 28568 31208 28580
rect 31260 28568 31266 28620
rect 37182 28608 37188 28620
rect 37143 28580 37188 28608
rect 37182 28568 37188 28580
rect 37240 28568 37246 28620
rect 46293 28611 46351 28617
rect 46293 28577 46305 28611
rect 46339 28608 46351 28611
rect 47026 28608 47032 28620
rect 46339 28580 47032 28608
rect 46339 28577 46351 28580
rect 46293 28571 46351 28577
rect 47026 28568 47032 28580
rect 47084 28568 47090 28620
rect 48130 28608 48136 28620
rect 48091 28580 48136 28608
rect 48130 28568 48136 28580
rect 48188 28568 48194 28620
rect 25455 28512 26096 28540
rect 26145 28543 26203 28549
rect 25455 28509 25467 28512
rect 25409 28503 25467 28509
rect 26145 28509 26157 28543
rect 26191 28509 26203 28543
rect 26145 28503 26203 28509
rect 17276 28444 18460 28472
rect 19696 28475 19754 28481
rect 17276 28432 17282 28444
rect 19696 28441 19708 28475
rect 19742 28472 19754 28475
rect 20070 28472 20076 28484
rect 19742 28444 20076 28472
rect 19742 28441 19754 28444
rect 19696 28435 19754 28441
rect 20070 28432 20076 28444
rect 20128 28432 20134 28484
rect 20180 28444 22094 28472
rect 12253 28407 12311 28413
rect 12253 28373 12265 28407
rect 12299 28404 12311 28407
rect 13081 28407 13139 28413
rect 13081 28404 13093 28407
rect 12299 28376 13093 28404
rect 12299 28373 12311 28376
rect 12253 28367 12311 28373
rect 13081 28373 13093 28376
rect 13127 28373 13139 28407
rect 13081 28367 13139 28373
rect 14093 28407 14151 28413
rect 14093 28373 14105 28407
rect 14139 28373 14151 28407
rect 14093 28367 14151 28373
rect 17678 28364 17684 28416
rect 17736 28404 17742 28416
rect 20180 28404 20208 28444
rect 20806 28404 20812 28416
rect 17736 28376 20208 28404
rect 20767 28376 20812 28404
rect 17736 28364 17742 28376
rect 20806 28364 20812 28376
rect 20864 28364 20870 28416
rect 22066 28404 22094 28444
rect 22278 28432 22284 28484
rect 22336 28472 22342 28484
rect 23658 28472 23664 28484
rect 22336 28444 23664 28472
rect 22336 28432 22342 28444
rect 23658 28432 23664 28444
rect 23716 28432 23722 28484
rect 24026 28432 24032 28484
rect 24084 28472 24090 28484
rect 26160 28472 26188 28503
rect 27982 28472 27988 28484
rect 24084 28444 26188 28472
rect 27943 28444 27988 28472
rect 24084 28432 24090 28444
rect 27982 28432 27988 28444
rect 28040 28432 28046 28484
rect 28169 28475 28227 28481
rect 28169 28441 28181 28475
rect 28215 28472 28227 28475
rect 29362 28472 29368 28484
rect 28215 28444 29368 28472
rect 28215 28441 28227 28444
rect 28169 28435 28227 28441
rect 29362 28432 29368 28444
rect 29420 28472 29426 28484
rect 30116 28472 30144 28568
rect 30834 28500 30840 28552
rect 30892 28540 30898 28552
rect 31461 28543 31519 28549
rect 31461 28540 31473 28543
rect 30892 28512 31473 28540
rect 30892 28500 30898 28512
rect 31461 28509 31473 28512
rect 31507 28509 31519 28543
rect 31461 28503 31519 28509
rect 32766 28500 32772 28552
rect 32824 28540 32830 28552
rect 33321 28543 33379 28549
rect 33321 28540 33333 28543
rect 32824 28512 33333 28540
rect 32824 28500 32830 28512
rect 33321 28509 33333 28512
rect 33367 28509 33379 28543
rect 33321 28503 33379 28509
rect 34606 28500 34612 28552
rect 34664 28540 34670 28552
rect 34701 28543 34759 28549
rect 34701 28540 34713 28543
rect 34664 28512 34713 28540
rect 34664 28500 34670 28512
rect 34701 28509 34713 28512
rect 34747 28509 34759 28543
rect 35526 28540 35532 28552
rect 35487 28512 35532 28540
rect 34701 28503 34759 28509
rect 35526 28500 35532 28512
rect 35584 28500 35590 28552
rect 29420 28444 30144 28472
rect 33873 28475 33931 28481
rect 29420 28432 29426 28444
rect 33873 28441 33885 28475
rect 33919 28472 33931 28475
rect 34054 28472 34060 28484
rect 33919 28444 34060 28472
rect 33919 28441 33931 28444
rect 33873 28435 33931 28441
rect 34054 28432 34060 28444
rect 34112 28432 34118 28484
rect 35710 28472 35716 28484
rect 35671 28444 35716 28472
rect 35710 28432 35716 28444
rect 35768 28432 35774 28484
rect 46477 28475 46535 28481
rect 46477 28441 46489 28475
rect 46523 28472 46535 28475
rect 47670 28472 47676 28484
rect 46523 28444 47676 28472
rect 46523 28441 46535 28444
rect 46477 28435 46535 28441
rect 47670 28432 47676 28444
rect 47728 28432 47734 28484
rect 24946 28404 24952 28416
rect 22066 28376 24952 28404
rect 24946 28364 24952 28376
rect 25004 28364 25010 28416
rect 25682 28404 25688 28416
rect 25643 28376 25688 28404
rect 25682 28364 25688 28376
rect 25740 28364 25746 28416
rect 28350 28404 28356 28416
rect 28311 28376 28356 28404
rect 28350 28364 28356 28376
rect 28408 28364 28414 28416
rect 32582 28404 32588 28416
rect 32543 28376 32588 28404
rect 32582 28364 32588 28376
rect 32640 28364 32646 28416
rect 1104 28314 48852 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 48852 28314
rect 1104 28240 48852 28262
rect 8018 28160 8024 28212
rect 8076 28200 8082 28212
rect 8076 28172 10732 28200
rect 8076 28160 8082 28172
rect 2866 28132 2872 28144
rect 2827 28104 2872 28132
rect 2866 28092 2872 28104
rect 2924 28092 2930 28144
rect 9852 28135 9910 28141
rect 7116 28104 8248 28132
rect 6914 28024 6920 28076
rect 6972 28064 6978 28076
rect 7116 28073 7144 28104
rect 8220 28076 8248 28104
rect 9852 28101 9864 28135
rect 9898 28132 9910 28135
rect 10594 28132 10600 28144
rect 9898 28104 10600 28132
rect 9898 28101 9910 28104
rect 9852 28095 9910 28101
rect 10594 28092 10600 28104
rect 10652 28092 10658 28144
rect 10704 28132 10732 28172
rect 12434 28160 12440 28212
rect 12492 28200 12498 28212
rect 12989 28203 13047 28209
rect 12989 28200 13001 28203
rect 12492 28172 13001 28200
rect 12492 28160 12498 28172
rect 12989 28169 13001 28172
rect 13035 28169 13047 28203
rect 12989 28163 13047 28169
rect 14274 28160 14280 28212
rect 14332 28200 14338 28212
rect 14369 28203 14427 28209
rect 14369 28200 14381 28203
rect 14332 28172 14381 28200
rect 14332 28160 14338 28172
rect 14369 28169 14381 28172
rect 14415 28169 14427 28203
rect 14369 28163 14427 28169
rect 16758 28160 16764 28212
rect 16816 28200 16822 28212
rect 17221 28203 17279 28209
rect 17221 28200 17233 28203
rect 16816 28172 17233 28200
rect 16816 28160 16822 28172
rect 17221 28169 17233 28172
rect 17267 28169 17279 28203
rect 17221 28163 17279 28169
rect 17957 28203 18015 28209
rect 17957 28169 17969 28203
rect 18003 28200 18015 28203
rect 19978 28200 19984 28212
rect 18003 28172 19984 28200
rect 18003 28169 18015 28172
rect 17957 28163 18015 28169
rect 19978 28160 19984 28172
rect 20036 28160 20042 28212
rect 23201 28203 23259 28209
rect 23201 28169 23213 28203
rect 23247 28200 23259 28203
rect 23566 28200 23572 28212
rect 23247 28172 23572 28200
rect 23247 28169 23259 28172
rect 23201 28163 23259 28169
rect 23566 28160 23572 28172
rect 23624 28160 23630 28212
rect 23658 28160 23664 28212
rect 23716 28200 23722 28212
rect 23716 28172 24624 28200
rect 23716 28160 23722 28172
rect 13814 28132 13820 28144
rect 10704 28104 12434 28132
rect 7101 28067 7159 28073
rect 7101 28064 7113 28067
rect 6972 28036 7113 28064
rect 6972 28024 6978 28036
rect 7101 28033 7113 28036
rect 7147 28033 7159 28067
rect 7101 28027 7159 28033
rect 7368 28067 7426 28073
rect 7368 28033 7380 28067
rect 7414 28064 7426 28067
rect 7414 28036 8156 28064
rect 7414 28033 7426 28036
rect 7368 28027 7426 28033
rect 2685 27999 2743 28005
rect 2685 27965 2697 27999
rect 2731 27965 2743 27999
rect 4154 27996 4160 28008
rect 4115 27968 4160 27996
rect 2685 27959 2743 27965
rect 2700 27928 2728 27959
rect 4154 27956 4160 27968
rect 4212 27956 4218 28008
rect 8128 27996 8156 28036
rect 8202 28024 8208 28076
rect 8260 28064 8266 28076
rect 9585 28067 9643 28073
rect 9585 28064 9597 28067
rect 8260 28036 9597 28064
rect 8260 28024 8266 28036
rect 9585 28033 9597 28036
rect 9631 28064 9643 28067
rect 9674 28064 9680 28076
rect 9631 28036 9680 28064
rect 9631 28033 9643 28036
rect 9585 28027 9643 28033
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 8938 27996 8944 28008
rect 8128 27968 8944 27996
rect 8938 27956 8944 27968
rect 8996 27956 9002 28008
rect 11238 27996 11244 28008
rect 10980 27968 11244 27996
rect 7006 27928 7012 27940
rect 2700 27900 7012 27928
rect 7006 27888 7012 27900
rect 7064 27888 7070 27940
rect 10980 27937 11008 27968
rect 11238 27956 11244 27968
rect 11296 27996 11302 28008
rect 11517 27999 11575 28005
rect 11517 27996 11529 27999
rect 11296 27968 11529 27996
rect 11296 27956 11302 27968
rect 11517 27965 11529 27968
rect 11563 27996 11575 27999
rect 11698 27996 11704 28008
rect 11563 27968 11704 27996
rect 11563 27965 11575 27968
rect 11517 27959 11575 27965
rect 11698 27956 11704 27968
rect 11756 27956 11762 28008
rect 11790 27956 11796 28008
rect 11848 27996 11854 28008
rect 12406 27996 12434 28104
rect 12912 28104 13820 28132
rect 12912 28073 12940 28104
rect 13814 28092 13820 28104
rect 13872 28132 13878 28144
rect 14001 28135 14059 28141
rect 14001 28132 14013 28135
rect 13872 28104 14013 28132
rect 13872 28092 13878 28104
rect 14001 28101 14013 28104
rect 14047 28101 14059 28135
rect 14001 28095 14059 28101
rect 14108 28104 15148 28132
rect 12897 28067 12955 28073
rect 12897 28033 12909 28067
rect 12943 28033 12955 28067
rect 12897 28027 12955 28033
rect 13081 28067 13139 28073
rect 13081 28033 13093 28067
rect 13127 28064 13139 28067
rect 14108 28064 14136 28104
rect 15120 28073 15148 28104
rect 18046 28092 18052 28144
rect 18104 28132 18110 28144
rect 19306 28135 19364 28141
rect 19306 28132 19318 28135
rect 18104 28104 19318 28132
rect 18104 28092 18110 28104
rect 19306 28101 19318 28104
rect 19352 28101 19364 28135
rect 24026 28132 24032 28144
rect 23987 28104 24032 28132
rect 19306 28095 19364 28101
rect 24026 28092 24032 28104
rect 24084 28092 24090 28144
rect 24596 28141 24624 28172
rect 25498 28160 25504 28212
rect 25556 28160 25562 28212
rect 27706 28160 27712 28212
rect 27764 28160 27770 28212
rect 35710 28160 35716 28212
rect 35768 28200 35774 28212
rect 37369 28203 37427 28209
rect 37369 28200 37381 28203
rect 35768 28172 37381 28200
rect 35768 28160 35774 28172
rect 37369 28169 37381 28172
rect 37415 28169 37427 28203
rect 37369 28163 37427 28169
rect 47670 28160 47676 28212
rect 47728 28200 47734 28212
rect 47854 28200 47860 28212
rect 47728 28172 47860 28200
rect 47728 28160 47734 28172
rect 47854 28160 47860 28172
rect 47912 28160 47918 28212
rect 24581 28135 24639 28141
rect 24581 28101 24593 28135
rect 24627 28101 24639 28135
rect 24581 28095 24639 28101
rect 24765 28135 24823 28141
rect 24765 28101 24777 28135
rect 24811 28132 24823 28135
rect 25130 28132 25136 28144
rect 24811 28104 25136 28132
rect 24811 28101 24823 28104
rect 24765 28095 24823 28101
rect 25130 28092 25136 28104
rect 25188 28092 25194 28144
rect 25516 28132 25544 28160
rect 25516 28104 25636 28132
rect 13127 28036 14136 28064
rect 14185 28067 14243 28073
rect 13127 28033 13139 28036
rect 13081 28027 13139 28033
rect 14185 28033 14197 28067
rect 14231 28033 14243 28067
rect 14185 28027 14243 28033
rect 15105 28067 15163 28073
rect 15105 28033 15117 28067
rect 15151 28064 15163 28067
rect 15838 28064 15844 28076
rect 15151 28036 15844 28064
rect 15151 28033 15163 28036
rect 15105 28027 15163 28033
rect 13096 27996 13124 28027
rect 11848 27968 11941 27996
rect 12406 27968 13124 27996
rect 14200 27996 14228 28027
rect 15838 28024 15844 28036
rect 15896 28024 15902 28076
rect 17126 28064 17132 28076
rect 17087 28036 17132 28064
rect 17126 28024 17132 28036
rect 17184 28024 17190 28076
rect 18230 28073 18236 28076
rect 18213 28067 18236 28073
rect 18213 28033 18225 28067
rect 18213 28027 18236 28033
rect 18230 28024 18236 28027
rect 18288 28024 18294 28076
rect 18322 28067 18380 28073
rect 18322 28033 18334 28067
rect 18368 28033 18380 28067
rect 18322 28027 18380 28033
rect 18417 28067 18475 28073
rect 18417 28033 18429 28067
rect 18463 28064 18475 28067
rect 18601 28067 18659 28073
rect 18463 28036 18552 28064
rect 18463 28033 18475 28036
rect 18417 28027 18475 28033
rect 14826 27996 14832 28008
rect 14200 27968 14832 27996
rect 11848 27956 11854 27968
rect 14826 27956 14832 27968
rect 14884 27956 14890 28008
rect 17218 27956 17224 28008
rect 17276 27996 17282 28008
rect 18337 27996 18365 28027
rect 17276 27968 18365 27996
rect 17276 27956 17282 27968
rect 10965 27931 11023 27937
rect 10965 27897 10977 27931
rect 11011 27897 11023 27931
rect 11808 27928 11836 27956
rect 17310 27928 17316 27940
rect 11808 27900 17316 27928
rect 10965 27891 11023 27897
rect 17310 27888 17316 27900
rect 17368 27888 17374 27940
rect 18524 27928 18552 28036
rect 18601 28033 18613 28067
rect 18647 28064 18659 28067
rect 19150 28064 19156 28076
rect 18647 28036 18736 28064
rect 18647 28033 18659 28036
rect 18601 28027 18659 28033
rect 18708 27996 18736 28036
rect 18984 28036 19156 28064
rect 18782 27996 18788 28008
rect 18708 27968 18788 27996
rect 18782 27956 18788 27968
rect 18840 27956 18846 28008
rect 18984 27928 19012 28036
rect 19150 28024 19156 28036
rect 19208 28024 19214 28076
rect 22465 28067 22523 28073
rect 22465 28033 22477 28067
rect 22511 28064 22523 28067
rect 23106 28064 23112 28076
rect 22511 28036 23112 28064
rect 22511 28033 22523 28036
rect 22465 28027 22523 28033
rect 23106 28024 23112 28036
rect 23164 28024 23170 28076
rect 25608 28073 25636 28104
rect 23845 28067 23903 28073
rect 23845 28033 23857 28067
rect 23891 28033 23903 28067
rect 23845 28027 23903 28033
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 25593 28067 25651 28073
rect 25593 28033 25605 28067
rect 25639 28033 25651 28067
rect 25593 28027 25651 28033
rect 19061 27999 19119 28005
rect 19061 27965 19073 27999
rect 19107 27965 19119 27999
rect 23860 27996 23888 28027
rect 24854 27996 24860 28008
rect 23860 27968 24860 27996
rect 19061 27959 19119 27965
rect 18524 27900 19012 27928
rect 8481 27863 8539 27869
rect 8481 27829 8493 27863
rect 8527 27860 8539 27863
rect 8570 27860 8576 27872
rect 8527 27832 8576 27860
rect 8527 27829 8539 27832
rect 8481 27823 8539 27829
rect 8570 27820 8576 27832
rect 8628 27820 8634 27872
rect 19076 27860 19104 27959
rect 24854 27956 24860 27968
rect 24912 27956 24918 28008
rect 25516 27996 25544 28027
rect 25682 28024 25688 28076
rect 25740 28064 25746 28076
rect 25740 28036 25785 28064
rect 25740 28024 25746 28036
rect 25866 28024 25872 28076
rect 25924 28064 25930 28076
rect 25924 28036 25969 28064
rect 25924 28024 25930 28036
rect 27430 28024 27436 28076
rect 27488 28064 27494 28076
rect 27724 28073 27752 28160
rect 29822 28132 29828 28144
rect 29380 28104 29828 28132
rect 27571 28067 27629 28073
rect 27571 28064 27583 28067
rect 27488 28036 27583 28064
rect 27488 28024 27494 28036
rect 27571 28033 27583 28036
rect 27617 28033 27629 28067
rect 27571 28027 27629 28033
rect 27709 28067 27767 28073
rect 27709 28033 27721 28067
rect 27755 28033 27767 28067
rect 27709 28027 27767 28033
rect 27806 28067 27864 28073
rect 27806 28033 27818 28067
rect 27852 28064 27864 28067
rect 27985 28067 28043 28073
rect 27852 28036 27936 28064
rect 27852 28033 27864 28036
rect 27806 28027 27864 28033
rect 26050 27996 26056 28008
rect 25516 27968 26056 27996
rect 26050 27956 26056 27968
rect 26108 27956 26114 28008
rect 27908 27996 27936 28036
rect 27985 28033 27997 28067
rect 28031 28064 28043 28067
rect 28350 28064 28356 28076
rect 28031 28036 28356 28064
rect 28031 28033 28043 28036
rect 27985 28027 28043 28033
rect 28350 28024 28356 28036
rect 28408 28024 28414 28076
rect 29270 28064 29276 28076
rect 29231 28036 29276 28064
rect 29270 28024 29276 28036
rect 29328 28024 29334 28076
rect 29380 28073 29408 28104
rect 29822 28092 29828 28104
rect 29880 28092 29886 28144
rect 34701 28135 34759 28141
rect 34701 28101 34713 28135
rect 34747 28132 34759 28135
rect 34790 28132 34796 28144
rect 34747 28104 34796 28132
rect 34747 28101 34759 28104
rect 34701 28095 34759 28101
rect 34790 28092 34796 28104
rect 34848 28092 34854 28144
rect 29365 28067 29423 28073
rect 29365 28033 29377 28067
rect 29411 28033 29423 28067
rect 29365 28027 29423 28033
rect 29457 28067 29515 28073
rect 29457 28033 29469 28067
rect 29503 28033 29515 28067
rect 29638 28064 29644 28076
rect 29599 28036 29644 28064
rect 29457 28027 29515 28033
rect 28902 27996 28908 28008
rect 27908 27968 28908 27996
rect 28902 27956 28908 27968
rect 28960 27996 28966 28008
rect 29472 27996 29500 28027
rect 29638 28024 29644 28036
rect 29696 28024 29702 28076
rect 30374 28024 30380 28076
rect 30432 28064 30438 28076
rect 30561 28067 30619 28073
rect 30561 28064 30573 28067
rect 30432 28036 30573 28064
rect 30432 28024 30438 28036
rect 30561 28033 30573 28036
rect 30607 28033 30619 28067
rect 32490 28064 32496 28076
rect 30561 28027 30619 28033
rect 30668 28036 32496 28064
rect 30668 27996 30696 28036
rect 32490 28024 32496 28036
rect 32548 28024 32554 28076
rect 32766 28064 32772 28076
rect 32727 28036 32772 28064
rect 32766 28024 32772 28036
rect 32824 28024 32830 28076
rect 33410 28024 33416 28076
rect 33468 28064 33474 28076
rect 34517 28067 34575 28073
rect 34517 28064 34529 28067
rect 33468 28036 34529 28064
rect 33468 28024 33474 28036
rect 34517 28033 34529 28036
rect 34563 28033 34575 28067
rect 37274 28064 37280 28076
rect 37235 28036 37280 28064
rect 34517 28027 34575 28033
rect 37274 28024 37280 28036
rect 37332 28024 37338 28076
rect 47854 28064 47860 28076
rect 47815 28036 47860 28064
rect 47854 28024 47860 28036
rect 47912 28024 47918 28076
rect 28960 27968 30696 27996
rect 28960 27956 28966 27968
rect 30742 27956 30748 28008
rect 30800 27996 30806 28008
rect 30929 27999 30987 28005
rect 30929 27996 30941 27999
rect 30800 27968 30941 27996
rect 30800 27956 30806 27968
rect 30929 27965 30941 27968
rect 30975 27996 30987 27999
rect 31294 27996 31300 28008
rect 30975 27968 31300 27996
rect 30975 27965 30987 27968
rect 30929 27959 30987 27965
rect 31294 27956 31300 27968
rect 31352 27956 31358 28008
rect 33226 27996 33232 28008
rect 33187 27968 33232 27996
rect 33226 27956 33232 27968
rect 33284 27956 33290 28008
rect 36357 27999 36415 28005
rect 36357 27965 36369 27999
rect 36403 27996 36415 27999
rect 36446 27996 36452 28008
rect 36403 27968 36452 27996
rect 36403 27965 36415 27968
rect 36357 27959 36415 27965
rect 36446 27956 36452 27968
rect 36504 27956 36510 28008
rect 27890 27888 27896 27940
rect 27948 27928 27954 27940
rect 35526 27928 35532 27940
rect 27948 27900 35532 27928
rect 27948 27888 27954 27900
rect 35526 27888 35532 27900
rect 35584 27888 35590 27940
rect 19426 27860 19432 27872
rect 19076 27832 19432 27860
rect 19426 27820 19432 27832
rect 19484 27860 19490 27872
rect 19702 27860 19708 27872
rect 19484 27832 19708 27860
rect 19484 27820 19490 27832
rect 19702 27820 19708 27832
rect 19760 27820 19766 27872
rect 20438 27860 20444 27872
rect 20399 27832 20444 27860
rect 20438 27820 20444 27832
rect 20496 27820 20502 27872
rect 22557 27863 22615 27869
rect 22557 27829 22569 27863
rect 22603 27860 22615 27863
rect 22738 27860 22744 27872
rect 22603 27832 22744 27860
rect 22603 27829 22615 27832
rect 22557 27823 22615 27829
rect 22738 27820 22744 27832
rect 22796 27820 22802 27872
rect 25225 27863 25283 27869
rect 25225 27829 25237 27863
rect 25271 27860 25283 27863
rect 25314 27860 25320 27872
rect 25271 27832 25320 27860
rect 25271 27829 25283 27832
rect 25225 27823 25283 27829
rect 25314 27820 25320 27832
rect 25372 27820 25378 27872
rect 27338 27860 27344 27872
rect 27299 27832 27344 27860
rect 27338 27820 27344 27832
rect 27396 27820 27402 27872
rect 28994 27860 29000 27872
rect 28955 27832 29000 27860
rect 28994 27820 29000 27832
rect 29052 27820 29058 27872
rect 48038 27860 48044 27872
rect 47999 27832 48044 27860
rect 48038 27820 48044 27832
rect 48096 27820 48102 27872
rect 1104 27770 48852 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 48852 27770
rect 1104 27696 48852 27718
rect 17218 27656 17224 27668
rect 10980 27628 11284 27656
rect 17179 27628 17224 27656
rect 8938 27588 8944 27600
rect 8899 27560 8944 27588
rect 8938 27548 8944 27560
rect 8996 27548 9002 27600
rect 10980 27588 11008 27628
rect 11256 27600 11284 27628
rect 17218 27616 17224 27628
rect 17276 27616 17282 27668
rect 20070 27656 20076 27668
rect 19352 27628 20076 27656
rect 11146 27588 11152 27600
rect 9048 27560 11008 27588
rect 11107 27560 11152 27588
rect 1394 27412 1400 27464
rect 1452 27452 1458 27464
rect 1581 27455 1639 27461
rect 1581 27452 1593 27455
rect 1452 27424 1593 27452
rect 1452 27412 1458 27424
rect 1581 27421 1593 27424
rect 1627 27421 1639 27455
rect 1581 27415 1639 27421
rect 2041 27455 2099 27461
rect 2041 27421 2053 27455
rect 2087 27452 2099 27455
rect 2222 27452 2228 27464
rect 2087 27424 2228 27452
rect 2087 27421 2099 27424
rect 2041 27415 2099 27421
rect 2222 27412 2228 27424
rect 2280 27412 2286 27464
rect 2869 27455 2927 27461
rect 2869 27452 2881 27455
rect 2746 27424 2881 27452
rect 1762 27344 1768 27396
rect 1820 27384 1826 27396
rect 2746 27384 2774 27424
rect 2869 27421 2881 27424
rect 2915 27421 2927 27455
rect 2869 27415 2927 27421
rect 6825 27455 6883 27461
rect 6825 27421 6837 27455
rect 6871 27452 6883 27455
rect 6914 27452 6920 27464
rect 6871 27424 6920 27452
rect 6871 27421 6883 27424
rect 6825 27415 6883 27421
rect 6914 27412 6920 27424
rect 6972 27412 6978 27464
rect 7092 27455 7150 27461
rect 7092 27421 7104 27455
rect 7138 27452 7150 27455
rect 8478 27452 8484 27464
rect 7138 27424 8484 27452
rect 7138 27421 7150 27424
rect 7092 27415 7150 27421
rect 8478 27412 8484 27424
rect 8536 27412 8542 27464
rect 1820 27356 2774 27384
rect 1820 27344 1826 27356
rect 3326 27344 3332 27396
rect 3384 27384 3390 27396
rect 9048 27384 9076 27560
rect 11146 27548 11152 27560
rect 11204 27548 11210 27600
rect 11238 27548 11244 27600
rect 11296 27548 11302 27600
rect 13078 27548 13084 27600
rect 13136 27588 13142 27600
rect 16114 27588 16120 27600
rect 13136 27560 16120 27588
rect 13136 27548 13142 27560
rect 16114 27548 16120 27560
rect 16172 27548 16178 27600
rect 16393 27591 16451 27597
rect 16393 27557 16405 27591
rect 16439 27588 16451 27591
rect 16666 27588 16672 27600
rect 16439 27560 16672 27588
rect 16439 27557 16451 27560
rect 16393 27551 16451 27557
rect 16666 27548 16672 27560
rect 16724 27548 16730 27600
rect 9122 27480 9128 27532
rect 9180 27520 9186 27532
rect 9180 27492 9444 27520
rect 9180 27480 9186 27492
rect 9416 27461 9444 27492
rect 9674 27480 9680 27532
rect 9732 27520 9738 27532
rect 11609 27523 11667 27529
rect 11609 27520 11621 27523
rect 9732 27492 11621 27520
rect 9732 27480 9738 27492
rect 11609 27489 11621 27492
rect 11655 27489 11667 27523
rect 11609 27483 11667 27489
rect 15746 27480 15752 27532
rect 15804 27520 15810 27532
rect 16574 27520 16580 27532
rect 15804 27492 16580 27520
rect 15804 27480 15810 27492
rect 16574 27480 16580 27492
rect 16632 27480 16638 27532
rect 17236 27520 17264 27616
rect 18049 27591 18107 27597
rect 18049 27557 18061 27591
rect 18095 27588 18107 27591
rect 19352 27588 19380 27628
rect 20070 27616 20076 27628
rect 20128 27616 20134 27668
rect 24946 27616 24952 27668
rect 25004 27656 25010 27668
rect 25682 27656 25688 27668
rect 25004 27628 25688 27656
rect 25004 27616 25010 27628
rect 25682 27616 25688 27628
rect 25740 27616 25746 27668
rect 27264 27628 28212 27656
rect 21082 27588 21088 27600
rect 18095 27560 19380 27588
rect 20995 27560 21088 27588
rect 18095 27557 18107 27560
rect 18049 27551 18107 27557
rect 21082 27548 21088 27560
rect 21140 27548 21146 27600
rect 22554 27548 22560 27600
rect 22612 27588 22618 27600
rect 27264 27588 27292 27628
rect 22612 27560 27292 27588
rect 28184 27588 28212 27628
rect 29564 27628 30512 27656
rect 29564 27588 29592 27628
rect 28184 27560 29592 27588
rect 30484 27588 30512 27628
rect 31680 27628 31800 27656
rect 31680 27588 31708 27628
rect 30484 27560 31708 27588
rect 31772 27588 31800 27628
rect 34606 27616 34612 27668
rect 34664 27656 34670 27668
rect 34885 27659 34943 27665
rect 34885 27656 34897 27659
rect 34664 27628 34897 27656
rect 34664 27616 34670 27628
rect 34885 27625 34897 27628
rect 34931 27625 34943 27659
rect 34885 27619 34943 27625
rect 33873 27591 33931 27597
rect 33873 27588 33885 27591
rect 31772 27560 33885 27588
rect 22612 27548 22618 27560
rect 33873 27557 33885 27560
rect 33919 27588 33931 27591
rect 34330 27588 34336 27600
rect 33919 27560 34336 27588
rect 33919 27557 33931 27560
rect 33873 27551 33931 27557
rect 34330 27548 34336 27560
rect 34388 27588 34394 27600
rect 47302 27588 47308 27600
rect 34388 27560 47308 27588
rect 34388 27548 34394 27560
rect 47302 27548 47308 27560
rect 47360 27548 47366 27600
rect 21100 27520 21128 27548
rect 25133 27523 25191 27529
rect 17236 27492 18460 27520
rect 21100 27492 21680 27520
rect 9217 27455 9275 27461
rect 9217 27421 9229 27455
rect 9263 27421 9275 27455
rect 9217 27415 9275 27421
rect 9309 27455 9367 27461
rect 9309 27421 9321 27455
rect 9355 27421 9367 27455
rect 9309 27415 9367 27421
rect 9401 27455 9459 27461
rect 9401 27421 9413 27455
rect 9447 27421 9459 27455
rect 9582 27452 9588 27464
rect 9543 27424 9588 27452
rect 9401 27415 9459 27421
rect 3384 27356 9076 27384
rect 3384 27344 3390 27356
rect 1946 27276 1952 27328
rect 2004 27316 2010 27328
rect 2133 27319 2191 27325
rect 2133 27316 2145 27319
rect 2004 27288 2145 27316
rect 2004 27276 2010 27288
rect 2133 27285 2145 27288
rect 2179 27285 2191 27319
rect 8202 27316 8208 27328
rect 8163 27288 8208 27316
rect 2133 27279 2191 27285
rect 8202 27276 8208 27288
rect 8260 27276 8266 27328
rect 9232 27316 9260 27415
rect 9324 27384 9352 27415
rect 9582 27412 9588 27424
rect 9640 27412 9646 27464
rect 11882 27461 11888 27464
rect 10137 27455 10195 27461
rect 10137 27421 10149 27455
rect 10183 27421 10195 27455
rect 10137 27415 10195 27421
rect 10321 27455 10379 27461
rect 10321 27421 10333 27455
rect 10367 27452 10379 27455
rect 11876 27452 11888 27461
rect 10367 27424 11008 27452
rect 11843 27424 11888 27452
rect 10367 27421 10379 27424
rect 10321 27415 10379 27421
rect 9490 27384 9496 27396
rect 9324 27356 9496 27384
rect 9490 27344 9496 27356
rect 9548 27344 9554 27396
rect 10152 27384 10180 27415
rect 10778 27384 10784 27396
rect 10152 27356 10784 27384
rect 10778 27344 10784 27356
rect 10836 27344 10842 27396
rect 10980 27393 11008 27424
rect 11876 27415 11888 27424
rect 11882 27412 11888 27415
rect 11940 27412 11946 27464
rect 16301 27455 16359 27461
rect 16301 27421 16313 27455
rect 16347 27452 16359 27455
rect 16390 27452 16396 27464
rect 16347 27424 16396 27452
rect 16347 27421 16359 27424
rect 16301 27415 16359 27421
rect 16390 27412 16396 27424
rect 16448 27412 16454 27464
rect 17126 27452 17132 27464
rect 16592 27424 17132 27452
rect 10965 27387 11023 27393
rect 10965 27353 10977 27387
rect 11011 27384 11023 27387
rect 11790 27384 11796 27396
rect 11011 27356 11796 27384
rect 11011 27353 11023 27356
rect 10965 27347 11023 27353
rect 11790 27344 11796 27356
rect 11848 27344 11854 27396
rect 16592 27393 16620 27424
rect 17126 27412 17132 27424
rect 17184 27412 17190 27464
rect 17310 27412 17316 27464
rect 17368 27452 17374 27464
rect 18432 27461 18460 27492
rect 18305 27455 18363 27461
rect 17368 27424 18276 27452
rect 17368 27412 17374 27424
rect 16577 27387 16635 27393
rect 12406 27356 16528 27384
rect 9766 27316 9772 27328
rect 9232 27288 9772 27316
rect 9766 27276 9772 27288
rect 9824 27316 9830 27328
rect 10226 27316 10232 27328
rect 9824 27288 10232 27316
rect 9824 27276 9830 27288
rect 10226 27276 10232 27288
rect 10284 27276 10290 27328
rect 10321 27319 10379 27325
rect 10321 27285 10333 27319
rect 10367 27316 10379 27319
rect 11054 27316 11060 27328
rect 10367 27288 11060 27316
rect 10367 27285 10379 27288
rect 10321 27279 10379 27285
rect 11054 27276 11060 27288
rect 11112 27276 11118 27328
rect 11238 27276 11244 27328
rect 11296 27316 11302 27328
rect 12406 27316 12434 27356
rect 11296 27288 12434 27316
rect 12989 27319 13047 27325
rect 11296 27276 11302 27288
rect 12989 27285 13001 27319
rect 13035 27316 13047 27319
rect 13262 27316 13268 27328
rect 13035 27288 13268 27316
rect 13035 27285 13047 27288
rect 12989 27279 13047 27285
rect 13262 27276 13268 27288
rect 13320 27276 13326 27328
rect 14274 27276 14280 27328
rect 14332 27316 14338 27328
rect 16298 27316 16304 27328
rect 14332 27288 16304 27316
rect 14332 27276 14338 27288
rect 16298 27276 16304 27288
rect 16356 27276 16362 27328
rect 16500 27316 16528 27356
rect 16577 27353 16589 27387
rect 16623 27353 16635 27387
rect 18248 27384 18276 27424
rect 18305 27421 18317 27455
rect 18351 27452 18363 27455
rect 18417 27455 18475 27461
rect 18351 27421 18368 27452
rect 18305 27415 18368 27421
rect 18417 27421 18429 27455
rect 18463 27421 18475 27455
rect 18530 27455 18588 27461
rect 18530 27452 18542 27455
rect 18417 27415 18475 27421
rect 18524 27421 18542 27452
rect 18576 27421 18588 27455
rect 18690 27452 18696 27464
rect 18651 27424 18696 27452
rect 18524 27415 18588 27421
rect 18340 27384 18368 27415
rect 16577 27347 16635 27353
rect 16684 27356 18184 27384
rect 18248 27356 18368 27384
rect 18524 27384 18552 27415
rect 18690 27412 18696 27424
rect 18748 27412 18754 27464
rect 19702 27452 19708 27464
rect 19663 27424 19708 27452
rect 19702 27412 19708 27424
rect 19760 27452 19766 27464
rect 21545 27455 21603 27461
rect 21545 27452 21557 27455
rect 19760 27424 21557 27452
rect 19760 27412 19766 27424
rect 21545 27421 21557 27424
rect 21591 27421 21603 27455
rect 21652 27452 21680 27492
rect 25133 27489 25145 27523
rect 25179 27520 25191 27523
rect 25774 27520 25780 27532
rect 25179 27492 25780 27520
rect 25179 27489 25191 27492
rect 25133 27483 25191 27489
rect 25774 27480 25780 27492
rect 25832 27480 25838 27532
rect 26786 27520 26792 27532
rect 26747 27492 26792 27520
rect 26786 27480 26792 27492
rect 26844 27480 26850 27532
rect 29546 27520 29552 27532
rect 29507 27492 29552 27520
rect 29546 27480 29552 27492
rect 29604 27480 29610 27532
rect 30558 27480 30564 27532
rect 30616 27520 30622 27532
rect 35621 27523 35679 27529
rect 35621 27520 35633 27523
rect 30616 27492 35633 27520
rect 30616 27480 30622 27492
rect 35621 27489 35633 27492
rect 35667 27489 35679 27523
rect 37090 27520 37096 27532
rect 37051 27492 37096 27520
rect 35621 27483 35679 27489
rect 37090 27480 37096 27492
rect 37148 27480 37154 27532
rect 23385 27455 23443 27461
rect 21652 27424 23336 27452
rect 21545 27415 21603 27421
rect 19334 27384 19340 27396
rect 18524 27356 19340 27384
rect 16684 27316 16712 27356
rect 16500 27288 16712 27316
rect 18156 27316 18184 27356
rect 19334 27344 19340 27356
rect 19392 27344 19398 27396
rect 19978 27393 19984 27396
rect 19972 27384 19984 27393
rect 19939 27356 19984 27384
rect 19972 27347 19984 27356
rect 19978 27344 19984 27347
rect 20036 27344 20042 27396
rect 20088 27356 21220 27384
rect 20088 27316 20116 27356
rect 18156 27288 20116 27316
rect 21192 27316 21220 27356
rect 21266 27344 21272 27396
rect 21324 27384 21330 27396
rect 21790 27387 21848 27393
rect 21790 27384 21802 27387
rect 21324 27356 21802 27384
rect 21324 27344 21330 27356
rect 21790 27353 21802 27356
rect 21836 27353 21848 27387
rect 23308 27384 23336 27424
rect 23385 27421 23397 27455
rect 23431 27452 23443 27455
rect 23658 27452 23664 27464
rect 23431 27424 23664 27452
rect 23431 27421 23443 27424
rect 23385 27415 23443 27421
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 24946 27452 24952 27464
rect 24907 27424 24952 27452
rect 24946 27412 24952 27424
rect 25004 27412 25010 27464
rect 27246 27452 27252 27464
rect 27207 27424 27252 27452
rect 27246 27412 27252 27424
rect 27304 27412 27310 27464
rect 27338 27412 27344 27464
rect 27396 27452 27402 27464
rect 27505 27455 27563 27461
rect 27505 27452 27517 27455
rect 27396 27424 27517 27452
rect 27396 27412 27402 27424
rect 27505 27421 27517 27424
rect 27551 27421 27563 27455
rect 27505 27415 27563 27421
rect 28994 27412 29000 27464
rect 29052 27452 29058 27464
rect 29805 27455 29863 27461
rect 29805 27452 29817 27455
rect 29052 27424 29817 27452
rect 29052 27412 29058 27424
rect 29805 27421 29817 27424
rect 29851 27421 29863 27455
rect 29805 27415 29863 27421
rect 31481 27455 31539 27461
rect 31481 27421 31493 27455
rect 31527 27452 31539 27455
rect 32401 27455 32459 27461
rect 32401 27452 32413 27455
rect 31527 27424 32413 27452
rect 31527 27421 31539 27424
rect 31481 27415 31539 27421
rect 32401 27421 32413 27424
rect 32447 27452 32459 27455
rect 32766 27452 32772 27464
rect 32447 27424 32772 27452
rect 32447 27421 32459 27424
rect 32401 27415 32459 27421
rect 32766 27412 32772 27424
rect 32824 27452 32830 27464
rect 34698 27452 34704 27464
rect 32824 27424 34704 27452
rect 32824 27412 32830 27424
rect 34698 27412 34704 27424
rect 34756 27412 34762 27464
rect 47302 27412 47308 27464
rect 47360 27452 47366 27464
rect 47670 27452 47676 27464
rect 47360 27424 47676 27452
rect 47360 27412 47366 27424
rect 47670 27412 47676 27424
rect 47728 27412 47734 27464
rect 31757 27387 31815 27393
rect 23308 27356 31064 27384
rect 21790 27347 21848 27353
rect 22462 27316 22468 27328
rect 21192 27288 22468 27316
rect 22462 27276 22468 27288
rect 22520 27276 22526 27328
rect 22554 27276 22560 27328
rect 22612 27316 22618 27328
rect 22925 27319 22983 27325
rect 22925 27316 22937 27319
rect 22612 27288 22937 27316
rect 22612 27276 22618 27288
rect 22925 27285 22937 27288
rect 22971 27285 22983 27319
rect 22925 27279 22983 27285
rect 23014 27276 23020 27328
rect 23072 27316 23078 27328
rect 23569 27319 23627 27325
rect 23569 27316 23581 27319
rect 23072 27288 23581 27316
rect 23072 27276 23078 27288
rect 23569 27285 23581 27288
rect 23615 27285 23627 27319
rect 28626 27316 28632 27328
rect 28587 27288 28632 27316
rect 23569 27279 23627 27285
rect 28626 27276 28632 27288
rect 28684 27276 28690 27328
rect 29178 27276 29184 27328
rect 29236 27316 29242 27328
rect 30929 27319 30987 27325
rect 30929 27316 30941 27319
rect 29236 27288 30941 27316
rect 29236 27276 29242 27288
rect 30929 27285 30941 27288
rect 30975 27285 30987 27319
rect 31036 27316 31064 27356
rect 31757 27353 31769 27387
rect 31803 27384 31815 27387
rect 33502 27384 33508 27396
rect 31803 27356 33508 27384
rect 31803 27353 31815 27356
rect 31757 27347 31815 27353
rect 33502 27344 33508 27356
rect 33560 27344 33566 27396
rect 35805 27387 35863 27393
rect 35805 27353 35817 27387
rect 35851 27384 35863 27387
rect 37366 27384 37372 27396
rect 35851 27356 37372 27384
rect 35851 27353 35863 27356
rect 35805 27347 35863 27353
rect 37366 27344 37372 27356
rect 37424 27344 37430 27396
rect 33594 27316 33600 27328
rect 31036 27288 33600 27316
rect 30929 27279 30987 27285
rect 33594 27276 33600 27288
rect 33652 27276 33658 27328
rect 1104 27226 48852 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 48852 27226
rect 1104 27152 48852 27174
rect 8481 27115 8539 27121
rect 8481 27081 8493 27115
rect 8527 27112 8539 27115
rect 9398 27112 9404 27124
rect 8527 27084 9404 27112
rect 8527 27081 8539 27084
rect 8481 27075 8539 27081
rect 9398 27072 9404 27084
rect 9456 27072 9462 27124
rect 9582 27072 9588 27124
rect 9640 27112 9646 27124
rect 13078 27112 13084 27124
rect 9640 27084 13084 27112
rect 9640 27072 9646 27084
rect 13078 27072 13084 27084
rect 13136 27072 13142 27124
rect 13262 27072 13268 27124
rect 13320 27112 13326 27124
rect 13541 27115 13599 27121
rect 13541 27112 13553 27115
rect 13320 27084 13553 27112
rect 13320 27072 13326 27084
rect 13541 27081 13553 27084
rect 13587 27081 13599 27115
rect 13541 27075 13599 27081
rect 13633 27115 13691 27121
rect 13633 27081 13645 27115
rect 13679 27112 13691 27115
rect 14366 27112 14372 27124
rect 13679 27084 14372 27112
rect 13679 27081 13691 27084
rect 13633 27075 13691 27081
rect 14366 27072 14372 27084
rect 14424 27072 14430 27124
rect 14826 27072 14832 27124
rect 14884 27112 14890 27124
rect 15010 27112 15016 27124
rect 14884 27084 15016 27112
rect 14884 27072 14890 27084
rect 15010 27072 15016 27084
rect 15068 27112 15074 27124
rect 15565 27115 15623 27121
rect 15565 27112 15577 27115
rect 15068 27084 15577 27112
rect 15068 27072 15074 27084
rect 15565 27081 15577 27084
rect 15611 27081 15623 27115
rect 15565 27075 15623 27081
rect 15654 27072 15660 27124
rect 15712 27112 15718 27124
rect 15712 27084 17816 27112
rect 15712 27072 15718 27084
rect 1946 27044 1952 27056
rect 1907 27016 1952 27044
rect 1946 27004 1952 27016
rect 2004 27004 2010 27056
rect 6546 27004 6552 27056
rect 6604 27044 6610 27056
rect 17313 27047 17371 27053
rect 6604 27016 16988 27044
rect 6604 27004 6610 27016
rect 1762 26976 1768 26988
rect 1723 26948 1768 26976
rect 1762 26936 1768 26948
rect 1820 26936 1826 26988
rect 7101 26979 7159 26985
rect 7101 26945 7113 26979
rect 7147 26976 7159 26979
rect 7190 26976 7196 26988
rect 7147 26948 7196 26976
rect 7147 26945 7159 26948
rect 7101 26939 7159 26945
rect 7190 26936 7196 26948
rect 7248 26936 7254 26988
rect 8018 26936 8024 26988
rect 8076 26976 8082 26988
rect 8113 26979 8171 26985
rect 8113 26976 8125 26979
rect 8076 26948 8125 26976
rect 8076 26936 8082 26948
rect 8113 26945 8125 26948
rect 8159 26945 8171 26979
rect 8113 26939 8171 26945
rect 8297 26979 8355 26985
rect 8297 26945 8309 26979
rect 8343 26945 8355 26979
rect 8297 26939 8355 26945
rect 2774 26868 2780 26920
rect 2832 26908 2838 26920
rect 2832 26880 2877 26908
rect 2832 26868 2838 26880
rect 7208 26840 7236 26936
rect 7374 26868 7380 26920
rect 7432 26908 7438 26920
rect 8202 26908 8208 26920
rect 7432 26880 8208 26908
rect 7432 26868 7438 26880
rect 8202 26868 8208 26880
rect 8260 26908 8266 26920
rect 8312 26908 8340 26939
rect 10778 26936 10784 26988
rect 10836 26976 10842 26988
rect 12618 26976 12624 26988
rect 10836 26948 12624 26976
rect 10836 26936 10842 26948
rect 12618 26936 12624 26948
rect 12676 26976 12682 26988
rect 13173 26979 13231 26985
rect 13173 26976 13185 26979
rect 12676 26948 13185 26976
rect 12676 26936 12682 26948
rect 13173 26945 13185 26948
rect 13219 26945 13231 26979
rect 13173 26939 13231 26945
rect 13449 26979 13507 26985
rect 13449 26945 13461 26979
rect 13495 26945 13507 26979
rect 13814 26976 13820 26988
rect 13775 26948 13820 26976
rect 13449 26939 13507 26945
rect 8260 26880 8340 26908
rect 13464 26908 13492 26939
rect 13814 26936 13820 26948
rect 13872 26936 13878 26988
rect 13909 26979 13967 26985
rect 13909 26945 13921 26979
rect 13955 26976 13967 26979
rect 15010 26976 15016 26988
rect 13955 26948 15016 26976
rect 13955 26945 13967 26948
rect 13909 26939 13967 26945
rect 15010 26936 15016 26948
rect 15068 26936 15074 26988
rect 15746 26976 15752 26988
rect 15707 26948 15752 26976
rect 15746 26936 15752 26948
rect 15804 26936 15810 26988
rect 15933 26979 15991 26985
rect 15933 26945 15945 26979
rect 15979 26976 15991 26979
rect 16666 26976 16672 26988
rect 15979 26948 16672 26976
rect 15979 26945 15991 26948
rect 15933 26939 15991 26945
rect 16666 26936 16672 26948
rect 16724 26936 16730 26988
rect 14090 26908 14096 26920
rect 13464 26880 14096 26908
rect 8260 26868 8266 26880
rect 14090 26868 14096 26880
rect 14148 26868 14154 26920
rect 14182 26868 14188 26920
rect 14240 26908 14246 26920
rect 14369 26911 14427 26917
rect 14369 26908 14381 26911
rect 14240 26880 14381 26908
rect 14240 26868 14246 26880
rect 14369 26877 14381 26880
rect 14415 26908 14427 26911
rect 15764 26908 15792 26936
rect 14415 26880 15792 26908
rect 16025 26911 16083 26917
rect 14415 26877 14427 26880
rect 14369 26871 14427 26877
rect 16025 26877 16037 26911
rect 16071 26908 16083 26911
rect 16390 26908 16396 26920
rect 16071 26880 16396 26908
rect 16071 26877 16083 26880
rect 16025 26871 16083 26877
rect 16390 26868 16396 26880
rect 16448 26868 16454 26920
rect 16960 26908 16988 27016
rect 17313 27013 17325 27047
rect 17359 27044 17371 27047
rect 17494 27044 17500 27056
rect 17359 27016 17500 27044
rect 17359 27013 17371 27016
rect 17313 27007 17371 27013
rect 17494 27004 17500 27016
rect 17552 27004 17558 27056
rect 17034 26936 17040 26988
rect 17092 26976 17098 26988
rect 17129 26979 17187 26985
rect 17129 26976 17141 26979
rect 17092 26948 17141 26976
rect 17092 26936 17098 26948
rect 17129 26945 17141 26948
rect 17175 26945 17187 26979
rect 17129 26939 17187 26945
rect 17402 26936 17408 26988
rect 17460 26976 17466 26988
rect 17788 26976 17816 27084
rect 18506 27072 18512 27124
rect 18564 27112 18570 27124
rect 19245 27115 19303 27121
rect 19245 27112 19257 27115
rect 18564 27084 19257 27112
rect 18564 27072 18570 27084
rect 19245 27081 19257 27084
rect 19291 27081 19303 27115
rect 19245 27075 19303 27081
rect 19334 27072 19340 27124
rect 19392 27112 19398 27124
rect 20073 27115 20131 27121
rect 20073 27112 20085 27115
rect 19392 27084 20085 27112
rect 19392 27072 19398 27084
rect 20073 27081 20085 27084
rect 20119 27081 20131 27115
rect 20073 27075 20131 27081
rect 20254 27072 20260 27124
rect 20312 27112 20318 27124
rect 24946 27112 24952 27124
rect 20312 27084 24952 27112
rect 20312 27072 20318 27084
rect 24946 27072 24952 27084
rect 25004 27072 25010 27124
rect 25038 27072 25044 27124
rect 25096 27112 25102 27124
rect 29549 27115 29607 27121
rect 25096 27084 29316 27112
rect 25096 27072 25102 27084
rect 17862 27004 17868 27056
rect 17920 27044 17926 27056
rect 18877 27047 18935 27053
rect 18877 27044 18889 27047
rect 17920 27016 18889 27044
rect 17920 27004 17926 27016
rect 18877 27013 18889 27016
rect 18923 27013 18935 27047
rect 18877 27007 18935 27013
rect 19061 27047 19119 27053
rect 19061 27013 19073 27047
rect 19107 27044 19119 27047
rect 19889 27047 19947 27053
rect 19107 27016 19840 27044
rect 19107 27013 19119 27016
rect 19061 27007 19119 27013
rect 18782 26976 18788 26988
rect 17460 26948 17505 26976
rect 17788 26948 18788 26976
rect 17460 26936 17466 26948
rect 18782 26936 18788 26948
rect 18840 26936 18846 26988
rect 18892 26976 18920 27007
rect 19705 26979 19763 26985
rect 19705 26976 19717 26979
rect 18892 26948 19717 26976
rect 19705 26945 19717 26948
rect 19751 26945 19763 26979
rect 19812 26976 19840 27016
rect 19889 27013 19901 27047
rect 19935 27044 19947 27047
rect 20806 27044 20812 27056
rect 19935 27016 20812 27044
rect 19935 27013 19947 27016
rect 19889 27007 19947 27013
rect 20806 27004 20812 27016
rect 20864 27004 20870 27056
rect 22738 27044 22744 27056
rect 22699 27016 22744 27044
rect 22738 27004 22744 27016
rect 22796 27004 22802 27056
rect 25314 27053 25320 27056
rect 25308 27007 25320 27053
rect 25372 27044 25378 27056
rect 27617 27047 27675 27053
rect 25372 27016 25408 27044
rect 25314 27004 25320 27007
rect 25372 27004 25378 27016
rect 27617 27013 27629 27047
rect 27663 27044 27675 27047
rect 28902 27044 28908 27056
rect 27663 27016 28908 27044
rect 27663 27013 27675 27016
rect 27617 27007 27675 27013
rect 28902 27004 28908 27016
rect 28960 27004 28966 27056
rect 29178 27044 29184 27056
rect 29139 27016 29184 27044
rect 29178 27004 29184 27016
rect 29236 27004 29242 27056
rect 29288 27044 29316 27084
rect 29549 27081 29561 27115
rect 29595 27112 29607 27115
rect 29638 27112 29644 27124
rect 29595 27084 29644 27112
rect 29595 27081 29607 27084
rect 29549 27075 29607 27081
rect 29638 27072 29644 27084
rect 29696 27072 29702 27124
rect 32122 27072 32128 27124
rect 32180 27112 32186 27124
rect 32493 27115 32551 27121
rect 32493 27112 32505 27115
rect 32180 27084 32505 27112
rect 32180 27072 32186 27084
rect 32493 27081 32505 27084
rect 32539 27081 32551 27115
rect 32493 27075 32551 27081
rect 34698 27072 34704 27124
rect 34756 27112 34762 27124
rect 35437 27115 35495 27121
rect 35437 27112 35449 27115
rect 34756 27084 35449 27112
rect 34756 27072 34762 27084
rect 35437 27081 35449 27084
rect 35483 27081 35495 27115
rect 35437 27075 35495 27081
rect 36173 27115 36231 27121
rect 36173 27081 36185 27115
rect 36219 27081 36231 27115
rect 37366 27112 37372 27124
rect 37327 27084 37372 27112
rect 36173 27075 36231 27081
rect 30558 27044 30564 27056
rect 29288 27016 30564 27044
rect 30558 27004 30564 27016
rect 30616 27004 30622 27056
rect 32309 27047 32367 27053
rect 32309 27013 32321 27047
rect 32355 27044 32367 27047
rect 32582 27044 32588 27056
rect 32355 27016 32588 27044
rect 32355 27013 32367 27016
rect 32309 27007 32367 27013
rect 32582 27004 32588 27016
rect 32640 27004 32646 27056
rect 33137 27047 33195 27053
rect 33137 27013 33149 27047
rect 33183 27044 33195 27047
rect 33686 27044 33692 27056
rect 33183 27016 33692 27044
rect 33183 27013 33195 27016
rect 33137 27007 33195 27013
rect 33686 27004 33692 27016
rect 33744 27004 33750 27056
rect 20438 26976 20444 26988
rect 19812 26948 20444 26976
rect 19705 26939 19763 26945
rect 20438 26936 20444 26948
rect 20496 26936 20502 26988
rect 22554 26976 22560 26988
rect 22515 26948 22560 26976
rect 22554 26936 22560 26948
rect 22612 26936 22618 26988
rect 25041 26979 25099 26985
rect 25041 26945 25053 26979
rect 25087 26976 25099 26979
rect 26326 26976 26332 26988
rect 25087 26974 25351 26976
rect 25424 26974 26332 26976
rect 25087 26948 26332 26974
rect 25087 26945 25099 26948
rect 25323 26946 25452 26948
rect 25041 26939 25099 26945
rect 26326 26936 26332 26948
rect 26384 26976 26390 26988
rect 27246 26976 27252 26988
rect 26384 26948 27252 26976
rect 26384 26936 26390 26948
rect 27246 26936 27252 26948
rect 27304 26936 27310 26988
rect 27430 26976 27436 26988
rect 27391 26948 27436 26976
rect 27430 26936 27436 26948
rect 27488 26936 27494 26988
rect 28166 26936 28172 26988
rect 28224 26976 28230 26988
rect 28537 26979 28595 26985
rect 28537 26976 28549 26979
rect 28224 26948 28549 26976
rect 28224 26936 28230 26948
rect 28537 26945 28549 26948
rect 28583 26945 28595 26979
rect 29362 26976 29368 26988
rect 29323 26948 29368 26976
rect 28537 26939 28595 26945
rect 29362 26936 29368 26948
rect 29420 26936 29426 26988
rect 30285 26979 30343 26985
rect 30285 26945 30297 26979
rect 30331 26976 30343 26979
rect 30374 26976 30380 26988
rect 30331 26948 30380 26976
rect 30331 26945 30343 26948
rect 30285 26939 30343 26945
rect 30374 26936 30380 26948
rect 30432 26936 30438 26988
rect 32125 26979 32183 26985
rect 32125 26945 32137 26979
rect 32171 26976 32183 26979
rect 32214 26976 32220 26988
rect 32171 26948 32220 26976
rect 32171 26945 32183 26948
rect 32125 26939 32183 26945
rect 32214 26936 32220 26948
rect 32272 26936 32278 26988
rect 32600 26976 32628 27004
rect 32953 26979 33011 26985
rect 32953 26976 32965 26979
rect 32600 26948 32965 26976
rect 32953 26945 32965 26948
rect 32999 26945 33011 26979
rect 34790 26976 34796 26988
rect 32953 26939 33011 26945
rect 34348 26948 34796 26976
rect 23750 26908 23756 26920
rect 16960 26880 18644 26908
rect 14274 26840 14280 26852
rect 7208 26812 14280 26840
rect 14274 26800 14280 26812
rect 14332 26800 14338 26852
rect 14737 26843 14795 26849
rect 14737 26809 14749 26843
rect 14783 26840 14795 26843
rect 15746 26840 15752 26852
rect 14783 26812 15752 26840
rect 14783 26809 14795 26812
rect 14737 26803 14795 26809
rect 15746 26800 15752 26812
rect 15804 26800 15810 26852
rect 16298 26800 16304 26852
rect 16356 26840 16362 26852
rect 18506 26840 18512 26852
rect 16356 26812 18512 26840
rect 16356 26800 16362 26812
rect 18506 26800 18512 26812
rect 18564 26800 18570 26852
rect 6730 26732 6736 26784
rect 6788 26772 6794 26784
rect 7193 26775 7251 26781
rect 7193 26772 7205 26775
rect 6788 26744 7205 26772
rect 6788 26732 6794 26744
rect 7193 26741 7205 26744
rect 7239 26741 7251 26775
rect 7193 26735 7251 26741
rect 13814 26732 13820 26784
rect 13872 26772 13878 26784
rect 14829 26775 14887 26781
rect 14829 26772 14841 26775
rect 13872 26744 14841 26772
rect 13872 26732 13878 26744
rect 14829 26741 14841 26744
rect 14875 26741 14887 26775
rect 14829 26735 14887 26741
rect 16758 26732 16764 26784
rect 16816 26772 16822 26784
rect 17129 26775 17187 26781
rect 17129 26772 17141 26775
rect 16816 26744 17141 26772
rect 16816 26732 16822 26744
rect 17129 26741 17141 26744
rect 17175 26741 17187 26775
rect 18616 26772 18644 26880
rect 18800 26880 23756 26908
rect 18800 26772 18828 26880
rect 23750 26868 23756 26880
rect 23808 26868 23814 26920
rect 23934 26908 23940 26920
rect 23895 26880 23940 26908
rect 23934 26868 23940 26880
rect 23992 26868 23998 26920
rect 26418 26868 26424 26920
rect 26476 26908 26482 26920
rect 26476 26880 30420 26908
rect 26476 26868 26482 26880
rect 18874 26800 18880 26852
rect 18932 26840 18938 26852
rect 19426 26840 19432 26852
rect 18932 26812 19432 26840
rect 18932 26800 18938 26812
rect 19426 26800 19432 26812
rect 19484 26840 19490 26852
rect 29546 26840 29552 26852
rect 19484 26812 25084 26840
rect 19484 26800 19490 26812
rect 18616 26744 18828 26772
rect 17129 26735 17187 26741
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 24946 26772 24952 26784
rect 20496 26744 24952 26772
rect 20496 26732 20502 26744
rect 24946 26732 24952 26744
rect 25004 26732 25010 26784
rect 25056 26772 25084 26812
rect 25976 26812 29552 26840
rect 25976 26772 26004 26812
rect 29546 26800 29552 26812
rect 29604 26800 29610 26852
rect 30392 26840 30420 26880
rect 30466 26868 30472 26920
rect 30524 26908 30530 26920
rect 30653 26911 30711 26917
rect 30653 26908 30665 26911
rect 30524 26880 30665 26908
rect 30524 26868 30530 26880
rect 30653 26877 30665 26880
rect 30699 26908 30711 26911
rect 31478 26908 31484 26920
rect 30699 26880 31484 26908
rect 30699 26877 30711 26880
rect 30653 26871 30711 26877
rect 31478 26868 31484 26880
rect 31536 26868 31542 26920
rect 32490 26868 32496 26920
rect 32548 26908 32554 26920
rect 34348 26908 34376 26948
rect 34790 26936 34796 26948
rect 34848 26976 34854 26988
rect 35253 26979 35311 26985
rect 35253 26976 35265 26979
rect 34848 26948 35265 26976
rect 34848 26936 34854 26948
rect 35253 26945 35265 26948
rect 35299 26945 35311 26979
rect 35253 26939 35311 26945
rect 35802 26936 35808 26988
rect 35860 26976 35866 26988
rect 35989 26979 36047 26985
rect 35989 26976 36001 26979
rect 35860 26948 36001 26976
rect 35860 26936 35866 26948
rect 35989 26945 36001 26948
rect 36035 26945 36047 26979
rect 36188 26976 36216 27075
rect 37366 27072 37372 27084
rect 37424 27072 37430 27124
rect 37274 26976 37280 26988
rect 36188 26948 37280 26976
rect 35989 26939 36047 26945
rect 37274 26936 37280 26948
rect 37332 26976 37338 26988
rect 37921 26979 37979 26985
rect 37921 26976 37933 26979
rect 37332 26948 37933 26976
rect 37332 26936 37338 26948
rect 37921 26945 37933 26948
rect 37967 26945 37979 26979
rect 37921 26939 37979 26945
rect 34698 26908 34704 26920
rect 32548 26880 34376 26908
rect 34659 26880 34704 26908
rect 32548 26868 32554 26880
rect 34698 26868 34704 26880
rect 34756 26868 34762 26920
rect 33318 26840 33324 26852
rect 30392 26812 33324 26840
rect 33318 26800 33324 26812
rect 33376 26800 33382 26852
rect 25056 26744 26004 26772
rect 26050 26732 26056 26784
rect 26108 26772 26114 26784
rect 26421 26775 26479 26781
rect 26421 26772 26433 26775
rect 26108 26744 26433 26772
rect 26108 26732 26114 26744
rect 26421 26741 26433 26744
rect 26467 26741 26479 26775
rect 26421 26735 26479 26741
rect 26694 26732 26700 26784
rect 26752 26772 26758 26784
rect 26878 26772 26884 26784
rect 26752 26744 26884 26772
rect 26752 26732 26758 26744
rect 26878 26732 26884 26744
rect 26936 26732 26942 26784
rect 27246 26732 27252 26784
rect 27304 26772 27310 26784
rect 27614 26772 27620 26784
rect 27304 26744 27620 26772
rect 27304 26732 27310 26744
rect 27614 26732 27620 26744
rect 27672 26732 27678 26784
rect 28629 26775 28687 26781
rect 28629 26741 28641 26775
rect 28675 26772 28687 26775
rect 29638 26772 29644 26784
rect 28675 26744 29644 26772
rect 28675 26741 28687 26744
rect 28629 26735 28687 26741
rect 29638 26732 29644 26744
rect 29696 26732 29702 26784
rect 36262 26732 36268 26784
rect 36320 26772 36326 26784
rect 38013 26775 38071 26781
rect 38013 26772 38025 26775
rect 36320 26744 38025 26772
rect 36320 26732 36326 26744
rect 38013 26741 38025 26744
rect 38059 26741 38071 26775
rect 38013 26735 38071 26741
rect 1104 26682 48852 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 48852 26682
rect 1104 26608 48852 26630
rect 3786 26528 3792 26580
rect 3844 26568 3850 26580
rect 15654 26568 15660 26580
rect 3844 26540 15660 26568
rect 3844 26528 3850 26540
rect 15654 26528 15660 26540
rect 15712 26528 15718 26580
rect 15746 26528 15752 26580
rect 15804 26568 15810 26580
rect 15804 26540 16620 26568
rect 15804 26528 15810 26540
rect 4798 26460 4804 26512
rect 4856 26500 4862 26512
rect 14734 26500 14740 26512
rect 4856 26472 7052 26500
rect 4856 26460 4862 26472
rect 1394 26432 1400 26444
rect 1355 26404 1400 26432
rect 1394 26392 1400 26404
rect 1452 26392 1458 26444
rect 2774 26392 2780 26444
rect 2832 26432 2838 26444
rect 6546 26432 6552 26444
rect 2832 26404 2877 26432
rect 6507 26404 6552 26432
rect 2832 26392 2838 26404
rect 6546 26392 6552 26404
rect 6604 26392 6610 26444
rect 6730 26432 6736 26444
rect 6691 26404 6736 26432
rect 6730 26392 6736 26404
rect 6788 26392 6794 26444
rect 7024 26441 7052 26472
rect 7944 26472 12434 26500
rect 14695 26472 14740 26500
rect 7009 26435 7067 26441
rect 7009 26401 7021 26435
rect 7055 26401 7067 26435
rect 7009 26395 7067 26401
rect 1578 26296 1584 26308
rect 1539 26268 1584 26296
rect 1578 26256 1584 26268
rect 1636 26256 1642 26308
rect 3970 26256 3976 26308
rect 4028 26296 4034 26308
rect 7944 26296 7972 26472
rect 8570 26392 8576 26444
rect 8628 26432 8634 26444
rect 8941 26435 8999 26441
rect 8941 26432 8953 26435
rect 8628 26404 8953 26432
rect 8628 26392 8634 26404
rect 8941 26401 8953 26404
rect 8987 26401 8999 26435
rect 10502 26432 10508 26444
rect 10463 26404 10508 26432
rect 8941 26395 8999 26401
rect 10502 26392 10508 26404
rect 10560 26392 10566 26444
rect 12406 26364 12434 26472
rect 14734 26460 14740 26472
rect 14792 26460 14798 26512
rect 16592 26432 16620 26540
rect 16666 26528 16672 26580
rect 16724 26568 16730 26580
rect 16761 26571 16819 26577
rect 16761 26568 16773 26571
rect 16724 26540 16773 26568
rect 16724 26528 16730 26540
rect 16761 26537 16773 26540
rect 16807 26568 16819 26571
rect 17034 26568 17040 26580
rect 16807 26540 17040 26568
rect 16807 26537 16819 26540
rect 16761 26531 16819 26537
rect 17034 26528 17040 26540
rect 17092 26568 17098 26580
rect 17221 26571 17279 26577
rect 17221 26568 17233 26571
rect 17092 26540 17233 26568
rect 17092 26528 17098 26540
rect 17221 26537 17233 26540
rect 17267 26537 17279 26571
rect 17221 26531 17279 26537
rect 17402 26528 17408 26580
rect 17460 26568 17466 26580
rect 18417 26571 18475 26577
rect 18417 26568 18429 26571
rect 17460 26540 18429 26568
rect 17460 26528 17466 26540
rect 18417 26537 18429 26540
rect 18463 26537 18475 26571
rect 18417 26531 18475 26537
rect 18506 26528 18512 26580
rect 18564 26568 18570 26580
rect 30834 26568 30840 26580
rect 18564 26540 30840 26568
rect 18564 26528 18570 26540
rect 30834 26528 30840 26540
rect 30892 26568 30898 26580
rect 46566 26568 46572 26580
rect 30892 26540 46572 26568
rect 30892 26528 30898 26540
rect 46566 26528 46572 26540
rect 46624 26528 46630 26580
rect 17494 26460 17500 26512
rect 17552 26500 17558 26512
rect 17589 26503 17647 26509
rect 17589 26500 17601 26503
rect 17552 26472 17601 26500
rect 17552 26460 17558 26472
rect 17589 26469 17601 26472
rect 17635 26469 17647 26503
rect 17589 26463 17647 26469
rect 17678 26460 17684 26512
rect 17736 26500 17742 26512
rect 24026 26500 24032 26512
rect 17736 26472 24032 26500
rect 17736 26460 17742 26472
rect 24026 26460 24032 26472
rect 24084 26460 24090 26512
rect 25133 26503 25191 26509
rect 25133 26469 25145 26503
rect 25179 26500 25191 26503
rect 25222 26500 25228 26512
rect 25179 26472 25228 26500
rect 25179 26469 25191 26472
rect 25133 26463 25191 26469
rect 25222 26460 25228 26472
rect 25280 26460 25286 26512
rect 25866 26460 25872 26512
rect 25924 26500 25930 26512
rect 45738 26500 45744 26512
rect 25924 26472 28994 26500
rect 25924 26460 25930 26472
rect 26050 26432 26056 26444
rect 16592 26404 18736 26432
rect 12406 26336 15332 26364
rect 9122 26296 9128 26308
rect 4028 26268 7972 26296
rect 9083 26268 9128 26296
rect 4028 26256 4034 26268
rect 9122 26256 9128 26268
rect 9180 26256 9186 26308
rect 13262 26256 13268 26308
rect 13320 26296 13326 26308
rect 14553 26299 14611 26305
rect 14553 26296 14565 26299
rect 13320 26268 14565 26296
rect 13320 26256 13326 26268
rect 14553 26265 14565 26268
rect 14599 26265 14611 26299
rect 15304 26296 15332 26336
rect 15378 26324 15384 26376
rect 15436 26364 15442 26376
rect 15436 26336 15481 26364
rect 15436 26324 15442 26336
rect 16390 26324 16396 26376
rect 16448 26364 16454 26376
rect 16448 26336 16804 26364
rect 16448 26324 16454 26336
rect 15470 26296 15476 26308
rect 15304 26268 15476 26296
rect 14553 26259 14611 26265
rect 15470 26256 15476 26268
rect 15528 26256 15534 26308
rect 15648 26299 15706 26305
rect 15648 26265 15660 26299
rect 15694 26296 15706 26299
rect 16666 26296 16672 26308
rect 15694 26268 16672 26296
rect 15694 26265 15706 26268
rect 15648 26259 15706 26265
rect 16666 26256 16672 26268
rect 16724 26256 16730 26308
rect 16776 26296 16804 26336
rect 17126 26324 17132 26376
rect 17184 26364 17190 26376
rect 17221 26367 17279 26373
rect 17221 26364 17233 26367
rect 17184 26336 17233 26364
rect 17184 26324 17190 26336
rect 17221 26333 17233 26336
rect 17267 26333 17279 26367
rect 17221 26327 17279 26333
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 18417 26367 18475 26373
rect 18417 26333 18429 26367
rect 18463 26364 18475 26367
rect 18598 26364 18604 26376
rect 18463 26336 18604 26364
rect 18463 26333 18475 26336
rect 18417 26327 18475 26333
rect 17420 26296 17448 26327
rect 18598 26324 18604 26336
rect 18656 26324 18662 26376
rect 18708 26373 18736 26404
rect 23492 26404 26056 26432
rect 18693 26367 18751 26373
rect 18693 26333 18705 26367
rect 18739 26364 18751 26367
rect 19426 26364 19432 26376
rect 18739 26336 19432 26364
rect 18739 26333 18751 26336
rect 18693 26327 18751 26333
rect 19426 26324 19432 26336
rect 19484 26324 19490 26376
rect 19521 26367 19579 26373
rect 19521 26333 19533 26367
rect 19567 26364 19579 26367
rect 20622 26364 20628 26376
rect 19567 26336 20628 26364
rect 19567 26333 19579 26336
rect 19521 26327 19579 26333
rect 20622 26324 20628 26336
rect 20680 26364 20686 26376
rect 23014 26364 23020 26376
rect 20680 26336 23020 26364
rect 20680 26324 20686 26336
rect 23014 26324 23020 26336
rect 23072 26324 23078 26376
rect 23492 26296 23520 26404
rect 26050 26392 26056 26404
rect 26108 26392 26114 26444
rect 26234 26392 26240 26444
rect 26292 26432 26298 26444
rect 27801 26435 27859 26441
rect 27801 26432 27813 26435
rect 26292 26404 27813 26432
rect 26292 26392 26298 26404
rect 27801 26401 27813 26404
rect 27847 26432 27859 26435
rect 28169 26435 28227 26441
rect 28169 26432 28181 26435
rect 27847 26404 28181 26432
rect 27847 26401 27859 26404
rect 27801 26395 27859 26401
rect 28169 26401 28181 26404
rect 28215 26401 28227 26435
rect 28169 26395 28227 26401
rect 26142 26364 26148 26376
rect 26103 26336 26148 26364
rect 26142 26324 26148 26336
rect 26200 26324 26206 26376
rect 27246 26364 27252 26376
rect 26252 26336 27252 26364
rect 23658 26296 23664 26308
rect 16776 26268 23520 26296
rect 23571 26268 23664 26296
rect 23658 26256 23664 26268
rect 23716 26296 23722 26308
rect 24762 26296 24768 26308
rect 23716 26268 24768 26296
rect 23716 26256 23722 26268
rect 24762 26256 24768 26268
rect 24820 26256 24826 26308
rect 24857 26299 24915 26305
rect 24857 26265 24869 26299
rect 24903 26296 24915 26299
rect 24946 26296 24952 26308
rect 24903 26268 24952 26296
rect 24903 26265 24915 26268
rect 24857 26259 24915 26265
rect 24946 26256 24952 26268
rect 25004 26256 25010 26308
rect 25682 26256 25688 26308
rect 25740 26296 25746 26308
rect 26252 26296 26280 26336
rect 27246 26324 27252 26336
rect 27304 26324 27310 26376
rect 27433 26367 27491 26373
rect 27433 26333 27445 26367
rect 27479 26364 27491 26367
rect 28276 26364 28304 26472
rect 28966 26432 28994 26472
rect 30576 26472 45744 26500
rect 30576 26432 30604 26472
rect 45738 26460 45744 26472
rect 45796 26460 45802 26512
rect 30834 26432 30840 26444
rect 28966 26404 30604 26432
rect 30795 26404 30840 26432
rect 30834 26392 30840 26404
rect 30892 26392 30898 26444
rect 32398 26432 32404 26444
rect 32359 26404 32404 26432
rect 32398 26392 32404 26404
rect 32456 26392 32462 26444
rect 33594 26392 33600 26444
rect 33652 26432 33658 26444
rect 35529 26435 35587 26441
rect 35529 26432 35541 26435
rect 33652 26404 35541 26432
rect 33652 26392 33658 26404
rect 35529 26401 35541 26404
rect 35575 26401 35587 26435
rect 35529 26395 35587 26401
rect 35713 26435 35771 26441
rect 35713 26401 35725 26435
rect 35759 26432 35771 26435
rect 36262 26432 36268 26444
rect 35759 26404 36268 26432
rect 35759 26401 35771 26404
rect 35713 26395 35771 26401
rect 36262 26392 36268 26404
rect 36320 26392 36326 26444
rect 45922 26432 45928 26444
rect 36924 26404 45928 26432
rect 28442 26364 28448 26376
rect 27479 26336 28304 26364
rect 28403 26336 28448 26364
rect 27479 26333 27491 26336
rect 27433 26327 27491 26333
rect 28442 26324 28448 26336
rect 28500 26324 28506 26376
rect 30193 26367 30251 26373
rect 30193 26333 30205 26367
rect 30239 26364 30251 26367
rect 31481 26367 31539 26373
rect 31481 26364 31493 26367
rect 30239 26336 31493 26364
rect 30239 26333 30251 26336
rect 30193 26327 30251 26333
rect 31481 26333 31493 26336
rect 31527 26364 31539 26367
rect 31938 26364 31944 26376
rect 31527 26336 31944 26364
rect 31527 26333 31539 26336
rect 31481 26327 31539 26333
rect 31938 26324 31944 26336
rect 31996 26324 32002 26376
rect 33505 26367 33563 26373
rect 33505 26364 33517 26367
rect 32416 26336 33517 26364
rect 25740 26268 26280 26296
rect 25740 26256 25746 26268
rect 26418 26256 26424 26308
rect 26476 26296 26482 26308
rect 26513 26299 26571 26305
rect 26513 26296 26525 26299
rect 26476 26268 26525 26296
rect 26476 26256 26482 26268
rect 26513 26265 26525 26268
rect 26559 26265 26571 26299
rect 26513 26259 26571 26265
rect 26620 26268 30328 26296
rect 2222 26188 2228 26240
rect 2280 26228 2286 26240
rect 17310 26228 17316 26240
rect 2280 26200 17316 26228
rect 2280 26188 2286 26200
rect 17310 26188 17316 26200
rect 17368 26188 17374 26240
rect 18230 26188 18236 26240
rect 18288 26228 18294 26240
rect 18601 26231 18659 26237
rect 18601 26228 18613 26231
rect 18288 26200 18613 26228
rect 18288 26188 18294 26200
rect 18601 26197 18613 26200
rect 18647 26228 18659 26231
rect 19242 26228 19248 26240
rect 18647 26200 19248 26228
rect 18647 26197 18659 26200
rect 18601 26191 18659 26197
rect 19242 26188 19248 26200
rect 19300 26188 19306 26240
rect 19705 26231 19763 26237
rect 19705 26197 19717 26231
rect 19751 26228 19763 26231
rect 20438 26228 20444 26240
rect 19751 26200 20444 26228
rect 19751 26197 19763 26200
rect 19705 26191 19763 26197
rect 20438 26188 20444 26200
rect 20496 26188 20502 26240
rect 23382 26188 23388 26240
rect 23440 26228 23446 26240
rect 23753 26231 23811 26237
rect 23753 26228 23765 26231
rect 23440 26200 23765 26228
rect 23440 26188 23446 26200
rect 23753 26197 23765 26200
rect 23799 26197 23811 26231
rect 23753 26191 23811 26197
rect 24026 26188 24032 26240
rect 24084 26228 24090 26240
rect 26620 26228 26648 26268
rect 27338 26228 27344 26240
rect 24084 26200 26648 26228
rect 27299 26200 27344 26228
rect 24084 26188 24090 26200
rect 27338 26188 27344 26200
rect 27396 26188 27402 26240
rect 30300 26228 30328 26268
rect 30374 26256 30380 26308
rect 30432 26296 30438 26308
rect 32416 26296 32444 26336
rect 33505 26333 33517 26336
rect 33551 26333 33563 26367
rect 33505 26327 33563 26333
rect 34701 26367 34759 26373
rect 34701 26333 34713 26367
rect 34747 26364 34759 26367
rect 34790 26364 34796 26376
rect 34747 26336 34796 26364
rect 34747 26333 34759 26336
rect 34701 26327 34759 26333
rect 30432 26268 32444 26296
rect 30432 26256 30438 26268
rect 30466 26228 30472 26240
rect 30300 26200 30472 26228
rect 30466 26188 30472 26200
rect 30524 26188 30530 26240
rect 33520 26228 33548 26327
rect 34790 26324 34796 26336
rect 34848 26324 34854 26376
rect 33962 26256 33968 26308
rect 34020 26296 34026 26308
rect 34057 26299 34115 26305
rect 34057 26296 34069 26299
rect 34020 26268 34069 26296
rect 34020 26256 34026 26268
rect 34057 26265 34069 26268
rect 34103 26296 34115 26299
rect 36924 26296 36952 26404
rect 45922 26392 45928 26404
rect 45980 26392 45986 26444
rect 34103 26268 36952 26296
rect 37369 26299 37427 26305
rect 34103 26265 34115 26268
rect 34057 26259 34115 26265
rect 37369 26265 37381 26299
rect 37415 26296 37427 26299
rect 44818 26296 44824 26308
rect 37415 26268 44824 26296
rect 37415 26265 37427 26268
rect 37369 26259 37427 26265
rect 44818 26256 44824 26268
rect 44876 26256 44882 26308
rect 47946 26296 47952 26308
rect 47907 26268 47952 26296
rect 47946 26256 47952 26268
rect 48004 26256 48010 26308
rect 48130 26296 48136 26308
rect 48091 26268 48136 26296
rect 48130 26256 48136 26268
rect 48188 26256 48194 26308
rect 34885 26231 34943 26237
rect 34885 26228 34897 26231
rect 33520 26200 34897 26228
rect 34885 26197 34897 26200
rect 34931 26228 34943 26231
rect 35158 26228 35164 26240
rect 34931 26200 35164 26228
rect 34931 26197 34943 26200
rect 34885 26191 34943 26197
rect 35158 26188 35164 26200
rect 35216 26228 35222 26240
rect 35802 26228 35808 26240
rect 35216 26200 35808 26228
rect 35216 26188 35222 26200
rect 35802 26188 35808 26200
rect 35860 26188 35866 26240
rect 1104 26138 48852 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 48852 26138
rect 1104 26064 48852 26086
rect 1578 25984 1584 26036
rect 1636 26024 1642 26036
rect 2317 26027 2375 26033
rect 2317 26024 2329 26027
rect 1636 25996 2329 26024
rect 1636 25984 1642 25996
rect 2317 25993 2329 25996
rect 2363 25993 2375 26027
rect 2317 25987 2375 25993
rect 2958 25984 2964 26036
rect 3016 26024 3022 26036
rect 8297 26027 8355 26033
rect 3016 25996 7420 26024
rect 3016 25984 3022 25996
rect 6365 25959 6423 25965
rect 6365 25925 6377 25959
rect 6411 25956 6423 25959
rect 6411 25928 7328 25956
rect 6411 25925 6423 25928
rect 6365 25919 6423 25925
rect 1578 25888 1584 25900
rect 1539 25860 1584 25888
rect 1578 25848 1584 25860
rect 1636 25848 1642 25900
rect 2222 25888 2228 25900
rect 2183 25860 2228 25888
rect 2222 25848 2228 25860
rect 2280 25848 2286 25900
rect 6638 25888 6644 25900
rect 6599 25860 6644 25888
rect 6638 25848 6644 25860
rect 6696 25848 6702 25900
rect 6270 25780 6276 25832
rect 6328 25820 6334 25832
rect 6457 25823 6515 25829
rect 6457 25820 6469 25823
rect 6328 25792 6469 25820
rect 6328 25780 6334 25792
rect 6457 25789 6469 25792
rect 6503 25789 6515 25823
rect 6457 25783 6515 25789
rect 1397 25755 1455 25761
rect 1397 25721 1409 25755
rect 1443 25752 1455 25755
rect 1443 25724 2774 25752
rect 1443 25721 1455 25724
rect 1397 25715 1455 25721
rect 2746 25684 2774 25724
rect 6365 25687 6423 25693
rect 6365 25684 6377 25687
rect 2746 25656 6377 25684
rect 6365 25653 6377 25656
rect 6411 25653 6423 25687
rect 6822 25684 6828 25696
rect 6783 25656 6828 25684
rect 6365 25647 6423 25653
rect 6822 25644 6828 25656
rect 6880 25644 6886 25696
rect 7300 25693 7328 25928
rect 7392 25752 7420 25996
rect 8297 25993 8309 26027
rect 8343 26024 8355 26027
rect 9122 26024 9128 26036
rect 8343 25996 9128 26024
rect 8343 25993 8355 25996
rect 8297 25987 8355 25993
rect 9122 25984 9128 25996
rect 9180 25984 9186 26036
rect 16666 26024 16672 26036
rect 16627 25996 16672 26024
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17034 26024 17040 26036
rect 16995 25996 17040 26024
rect 17034 25984 17040 25996
rect 17092 25984 17098 26036
rect 25222 26024 25228 26036
rect 17236 25996 25228 26024
rect 17236 25956 17264 25996
rect 25222 25984 25228 25996
rect 25280 25984 25286 26036
rect 28166 26024 28172 26036
rect 26252 25996 28172 26024
rect 8220 25928 17264 25956
rect 7742 25848 7748 25900
rect 7800 25888 7806 25900
rect 8220 25897 8248 25928
rect 17402 25916 17408 25968
rect 17460 25956 17466 25968
rect 26050 25956 26056 25968
rect 17460 25928 26056 25956
rect 17460 25916 17466 25928
rect 26050 25916 26056 25928
rect 26108 25956 26114 25968
rect 26252 25965 26280 25996
rect 28166 25984 28172 25996
rect 28224 25984 28230 26036
rect 28442 25984 28448 26036
rect 28500 26024 28506 26036
rect 28500 25996 31754 26024
rect 28500 25984 28506 25996
rect 26237 25959 26295 25965
rect 26237 25956 26249 25959
rect 26108 25928 26249 25956
rect 26108 25916 26114 25928
rect 26237 25925 26249 25928
rect 26283 25925 26295 25959
rect 26237 25919 26295 25925
rect 26970 25916 26976 25968
rect 27028 25956 27034 25968
rect 28261 25959 28319 25965
rect 28261 25956 28273 25959
rect 27028 25928 28273 25956
rect 27028 25916 27034 25928
rect 28261 25925 28273 25928
rect 28307 25956 28319 25959
rect 28350 25956 28356 25968
rect 28307 25928 28356 25956
rect 28307 25925 28319 25928
rect 28261 25919 28319 25925
rect 28350 25916 28356 25928
rect 28408 25916 28414 25968
rect 8205 25891 8263 25897
rect 8205 25888 8217 25891
rect 7800 25860 8217 25888
rect 7800 25848 7806 25860
rect 8205 25857 8217 25860
rect 8251 25857 8263 25891
rect 8205 25851 8263 25857
rect 8294 25848 8300 25900
rect 8352 25888 8358 25900
rect 9306 25888 9312 25900
rect 8352 25860 9312 25888
rect 8352 25848 8358 25860
rect 9306 25848 9312 25860
rect 9364 25848 9370 25900
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 11701 25891 11759 25897
rect 11701 25888 11713 25891
rect 10284 25860 11713 25888
rect 10284 25848 10290 25860
rect 11701 25857 11713 25860
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 13081 25891 13139 25897
rect 13081 25857 13093 25891
rect 13127 25857 13139 25891
rect 13262 25888 13268 25900
rect 13223 25860 13268 25888
rect 13081 25851 13139 25857
rect 9214 25780 9220 25832
rect 9272 25820 9278 25832
rect 9585 25823 9643 25829
rect 9585 25820 9597 25823
rect 9272 25792 9597 25820
rect 9272 25780 9278 25792
rect 9585 25789 9597 25792
rect 9631 25789 9643 25823
rect 11606 25820 11612 25832
rect 11567 25792 11612 25820
rect 9585 25783 9643 25789
rect 11606 25780 11612 25792
rect 11664 25780 11670 25832
rect 13096 25820 13124 25851
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 14182 25888 14188 25900
rect 14143 25860 14188 25888
rect 14182 25848 14188 25860
rect 14240 25848 14246 25900
rect 16853 25891 16911 25897
rect 16853 25857 16865 25891
rect 16899 25886 16911 25891
rect 16942 25886 16948 25900
rect 16899 25858 16948 25886
rect 16899 25857 16911 25858
rect 16853 25851 16911 25857
rect 16942 25848 16948 25858
rect 17000 25848 17006 25900
rect 17126 25888 17132 25900
rect 17087 25860 17132 25888
rect 17126 25848 17132 25860
rect 17184 25848 17190 25900
rect 18500 25891 18558 25897
rect 18500 25857 18512 25891
rect 18546 25888 18558 25891
rect 20257 25891 20315 25897
rect 20257 25888 20269 25891
rect 18546 25860 20269 25888
rect 18546 25857 18558 25860
rect 18500 25851 18558 25857
rect 20257 25857 20269 25860
rect 20303 25857 20315 25891
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20257 25851 20315 25857
rect 20364 25860 20453 25888
rect 14274 25820 14280 25832
rect 13096 25792 14280 25820
rect 14274 25780 14280 25792
rect 14332 25780 14338 25832
rect 18230 25820 18236 25832
rect 18191 25792 18236 25820
rect 18230 25780 18236 25792
rect 18288 25780 18294 25832
rect 19518 25780 19524 25832
rect 19576 25820 19582 25832
rect 20073 25823 20131 25829
rect 20073 25820 20085 25823
rect 19576 25792 20085 25820
rect 19576 25780 19582 25792
rect 20073 25789 20085 25792
rect 20119 25789 20131 25823
rect 20073 25783 20131 25789
rect 12710 25752 12716 25764
rect 7392 25724 12716 25752
rect 12710 25712 12716 25724
rect 12768 25712 12774 25764
rect 19242 25712 19248 25764
rect 19300 25752 19306 25764
rect 20364 25752 20392 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20533 25891 20591 25897
rect 20533 25857 20545 25891
rect 20579 25857 20591 25891
rect 23474 25888 23480 25900
rect 23435 25860 23480 25888
rect 20533 25851 20591 25857
rect 20548 25820 20576 25851
rect 23474 25848 23480 25860
rect 23532 25848 23538 25900
rect 23753 25891 23811 25897
rect 23753 25857 23765 25891
rect 23799 25857 23811 25891
rect 24578 25888 24584 25900
rect 24491 25860 24584 25888
rect 23753 25851 23811 25857
rect 23566 25820 23572 25832
rect 20456 25792 20576 25820
rect 23527 25792 23572 25820
rect 20456 25764 20484 25792
rect 23566 25780 23572 25792
rect 23624 25780 23630 25832
rect 23768 25820 23796 25851
rect 24578 25848 24584 25860
rect 24636 25888 24642 25900
rect 25777 25891 25835 25897
rect 25777 25888 25789 25891
rect 24636 25860 25789 25888
rect 24636 25848 24642 25860
rect 25777 25857 25789 25860
rect 25823 25888 25835 25891
rect 26142 25888 26148 25900
rect 25823 25860 26148 25888
rect 25823 25857 25835 25860
rect 25777 25851 25835 25857
rect 26142 25848 26148 25860
rect 26200 25848 26206 25900
rect 27065 25891 27123 25897
rect 27065 25857 27077 25891
rect 27111 25888 27123 25891
rect 27893 25891 27951 25897
rect 27893 25888 27905 25891
rect 27111 25860 27905 25888
rect 27111 25857 27123 25860
rect 27065 25851 27123 25857
rect 27893 25857 27905 25860
rect 27939 25888 27951 25891
rect 28460 25888 28488 25984
rect 29638 25956 29644 25968
rect 29599 25928 29644 25956
rect 29638 25916 29644 25928
rect 29696 25916 29702 25968
rect 27939 25860 28488 25888
rect 27939 25857 27951 25860
rect 27893 25851 27951 25857
rect 29178 25848 29184 25900
rect 29236 25888 29242 25900
rect 29457 25891 29515 25897
rect 29457 25888 29469 25891
rect 29236 25860 29469 25888
rect 29236 25848 29242 25860
rect 29457 25857 29469 25860
rect 29503 25857 29515 25891
rect 31726 25888 31754 25996
rect 32030 25916 32036 25968
rect 32088 25956 32094 25968
rect 34701 25959 34759 25965
rect 32088 25928 34284 25956
rect 32088 25916 32094 25928
rect 32125 25891 32183 25897
rect 32125 25888 32137 25891
rect 31726 25860 32137 25888
rect 29457 25851 29515 25857
rect 32125 25857 32137 25860
rect 32171 25888 32183 25891
rect 32490 25888 32496 25900
rect 32171 25860 32496 25888
rect 32171 25857 32183 25860
rect 32125 25851 32183 25857
rect 32490 25848 32496 25860
rect 32548 25848 32554 25900
rect 23768 25792 25084 25820
rect 19300 25724 20392 25752
rect 19300 25712 19306 25724
rect 20438 25712 20444 25764
rect 20496 25712 20502 25764
rect 22370 25712 22376 25764
rect 22428 25752 22434 25764
rect 24854 25752 24860 25764
rect 22428 25724 24860 25752
rect 22428 25712 22434 25724
rect 24854 25712 24860 25724
rect 24912 25712 24918 25764
rect 7285 25687 7343 25693
rect 7285 25653 7297 25687
rect 7331 25684 7343 25687
rect 10962 25684 10968 25696
rect 7331 25656 10968 25684
rect 7331 25653 7343 25656
rect 7285 25647 7343 25653
rect 10962 25644 10968 25656
rect 11020 25644 11026 25696
rect 11977 25687 12035 25693
rect 11977 25653 11989 25687
rect 12023 25684 12035 25687
rect 12066 25684 12072 25696
rect 12023 25656 12072 25684
rect 12023 25653 12035 25656
rect 11977 25647 12035 25653
rect 12066 25644 12072 25656
rect 12124 25644 12130 25696
rect 12250 25644 12256 25696
rect 12308 25684 12314 25696
rect 13173 25687 13231 25693
rect 13173 25684 13185 25687
rect 12308 25656 13185 25684
rect 12308 25644 12314 25656
rect 13173 25653 13185 25656
rect 13219 25653 13231 25687
rect 13173 25647 13231 25653
rect 16942 25644 16948 25696
rect 17000 25684 17006 25696
rect 17402 25684 17408 25696
rect 17000 25656 17408 25684
rect 17000 25644 17006 25656
rect 17402 25644 17408 25656
rect 17460 25644 17466 25696
rect 18230 25644 18236 25696
rect 18288 25684 18294 25696
rect 19426 25684 19432 25696
rect 18288 25656 19432 25684
rect 18288 25644 18294 25656
rect 19426 25644 19432 25656
rect 19484 25644 19490 25696
rect 19610 25684 19616 25696
rect 19571 25656 19616 25684
rect 19610 25644 19616 25656
rect 19668 25644 19674 25696
rect 19702 25644 19708 25696
rect 19760 25684 19766 25696
rect 23477 25687 23535 25693
rect 23477 25684 23489 25687
rect 19760 25656 23489 25684
rect 19760 25644 19766 25656
rect 23477 25653 23489 25656
rect 23523 25653 23535 25687
rect 23934 25684 23940 25696
rect 23895 25656 23940 25684
rect 23477 25647 23535 25653
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 25056 25684 25084 25792
rect 25130 25780 25136 25832
rect 25188 25820 25194 25832
rect 25498 25820 25504 25832
rect 25188 25792 25504 25820
rect 25188 25780 25194 25792
rect 25498 25780 25504 25792
rect 25556 25780 25562 25832
rect 31018 25820 31024 25832
rect 30979 25792 31024 25820
rect 31018 25780 31024 25792
rect 31076 25780 31082 25832
rect 31570 25780 31576 25832
rect 31628 25820 31634 25832
rect 32861 25823 32919 25829
rect 32861 25820 32873 25823
rect 31628 25792 32873 25820
rect 31628 25780 31634 25792
rect 32861 25789 32873 25792
rect 32907 25789 32919 25823
rect 33042 25820 33048 25832
rect 33003 25792 33048 25820
rect 32861 25783 32919 25789
rect 33042 25780 33048 25792
rect 33100 25780 33106 25832
rect 34256 25820 34284 25928
rect 34701 25925 34713 25959
rect 34747 25956 34759 25959
rect 45554 25956 45560 25968
rect 34747 25928 45560 25956
rect 34747 25925 34759 25928
rect 34701 25919 34759 25925
rect 45554 25916 45560 25928
rect 45612 25916 45618 25968
rect 35158 25888 35164 25900
rect 35119 25860 35164 25888
rect 35158 25848 35164 25860
rect 35216 25848 35222 25900
rect 35802 25820 35808 25832
rect 34256 25792 35808 25820
rect 35802 25780 35808 25792
rect 35860 25820 35866 25832
rect 46658 25820 46664 25832
rect 35860 25792 46664 25820
rect 35860 25780 35866 25792
rect 46658 25780 46664 25792
rect 46716 25780 46722 25832
rect 25222 25712 25228 25764
rect 25280 25752 25286 25764
rect 33962 25752 33968 25764
rect 25280 25724 33968 25752
rect 25280 25712 25286 25724
rect 33962 25712 33968 25724
rect 34020 25712 34026 25764
rect 27154 25684 27160 25696
rect 25056 25656 27160 25684
rect 27154 25644 27160 25656
rect 27212 25644 27218 25696
rect 27249 25687 27307 25693
rect 27249 25653 27261 25687
rect 27295 25684 27307 25687
rect 27982 25684 27988 25696
rect 27295 25656 27988 25684
rect 27295 25653 27307 25656
rect 27249 25647 27307 25653
rect 27982 25644 27988 25656
rect 28040 25644 28046 25696
rect 31938 25644 31944 25696
rect 31996 25684 32002 25696
rect 32309 25687 32367 25693
rect 32309 25684 32321 25687
rect 31996 25656 32321 25684
rect 31996 25644 32002 25656
rect 32309 25653 32321 25656
rect 32355 25684 32367 25687
rect 32490 25684 32496 25696
rect 32355 25656 32496 25684
rect 32355 25653 32367 25656
rect 32309 25647 32367 25653
rect 32490 25644 32496 25656
rect 32548 25644 32554 25696
rect 1104 25594 48852 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 48852 25594
rect 1104 25520 48852 25542
rect 6822 25440 6828 25492
rect 6880 25480 6886 25492
rect 19702 25480 19708 25492
rect 6880 25452 19708 25480
rect 6880 25440 6886 25452
rect 19702 25440 19708 25452
rect 19760 25440 19766 25492
rect 23198 25480 23204 25492
rect 20548 25452 21487 25480
rect 23159 25452 23204 25480
rect 8128 25384 9444 25412
rect 8128 25285 8156 25384
rect 9214 25344 9220 25356
rect 9175 25316 9220 25344
rect 9214 25304 9220 25316
rect 9272 25304 9278 25356
rect 9416 25344 9444 25384
rect 9766 25372 9772 25424
rect 9824 25412 9830 25424
rect 10778 25412 10784 25424
rect 9824 25384 10784 25412
rect 9824 25372 9830 25384
rect 10778 25372 10784 25384
rect 10836 25372 10842 25424
rect 11330 25372 11336 25424
rect 11388 25412 11394 25424
rect 11793 25415 11851 25421
rect 11793 25412 11805 25415
rect 11388 25384 11805 25412
rect 11388 25372 11394 25384
rect 11793 25381 11805 25384
rect 11839 25381 11851 25415
rect 12066 25412 12072 25424
rect 12027 25384 12072 25412
rect 11793 25375 11851 25381
rect 12066 25372 12072 25384
rect 12124 25372 12130 25424
rect 13170 25372 13176 25424
rect 13228 25412 13234 25424
rect 14458 25412 14464 25424
rect 13228 25384 14464 25412
rect 13228 25372 13234 25384
rect 9677 25347 9735 25353
rect 9677 25344 9689 25347
rect 9416 25316 9689 25344
rect 9677 25313 9689 25316
rect 9723 25344 9735 25347
rect 9858 25344 9864 25356
rect 9723 25316 9864 25344
rect 9723 25313 9735 25316
rect 9677 25307 9735 25313
rect 9858 25304 9864 25316
rect 9916 25304 9922 25356
rect 10321 25347 10379 25353
rect 10321 25313 10333 25347
rect 10367 25344 10379 25347
rect 12161 25347 12219 25353
rect 10367 25316 12020 25344
rect 10367 25313 10379 25316
rect 10321 25307 10379 25313
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 8113 25279 8171 25285
rect 8113 25245 8125 25279
rect 8159 25245 8171 25279
rect 8113 25239 8171 25245
rect 8205 25279 8263 25285
rect 8205 25245 8217 25279
rect 8251 25276 8263 25279
rect 8754 25276 8760 25288
rect 8251 25248 8760 25276
rect 8251 25245 8263 25248
rect 8205 25239 8263 25245
rect 8036 25208 8064 25239
rect 8754 25236 8760 25248
rect 8812 25276 8818 25288
rect 9582 25276 9588 25288
rect 8812 25248 9588 25276
rect 8812 25236 8818 25248
rect 9582 25236 9588 25248
rect 9640 25236 9646 25288
rect 10505 25279 10563 25285
rect 10505 25276 10517 25279
rect 9784 25248 10517 25276
rect 8294 25208 8300 25220
rect 8036 25180 8300 25208
rect 8294 25168 8300 25180
rect 8352 25168 8358 25220
rect 8389 25211 8447 25217
rect 8389 25177 8401 25211
rect 8435 25208 8447 25211
rect 9784 25208 9812 25248
rect 10505 25245 10517 25248
rect 10551 25245 10563 25279
rect 10505 25239 10563 25245
rect 10597 25279 10655 25285
rect 10597 25245 10609 25279
rect 10643 25245 10655 25279
rect 10778 25276 10784 25288
rect 10739 25248 10784 25276
rect 10597 25239 10655 25245
rect 8435 25180 9812 25208
rect 9861 25211 9919 25217
rect 8435 25177 8447 25180
rect 8389 25171 8447 25177
rect 9861 25177 9873 25211
rect 9907 25208 9919 25211
rect 10612 25208 10640 25239
rect 10778 25236 10784 25248
rect 10836 25236 10842 25288
rect 10870 25236 10876 25288
rect 10928 25276 10934 25288
rect 11992 25285 12020 25316
rect 12161 25313 12173 25347
rect 12207 25344 12219 25347
rect 12986 25344 12992 25356
rect 12207 25316 12992 25344
rect 12207 25313 12219 25316
rect 12161 25307 12219 25313
rect 12986 25304 12992 25316
rect 13044 25304 13050 25356
rect 13280 25353 13308 25384
rect 14458 25372 14464 25384
rect 14516 25372 14522 25424
rect 17310 25372 17316 25424
rect 17368 25412 17374 25424
rect 20548 25412 20576 25452
rect 17368 25384 20576 25412
rect 21459 25412 21487 25452
rect 23198 25440 23204 25452
rect 23256 25440 23262 25492
rect 23566 25480 23572 25492
rect 23527 25452 23572 25480
rect 23566 25440 23572 25452
rect 23624 25440 23630 25492
rect 25130 25480 25136 25492
rect 23676 25452 25136 25480
rect 23676 25412 23704 25452
rect 25130 25440 25136 25452
rect 25188 25440 25194 25492
rect 25501 25483 25559 25489
rect 25501 25449 25513 25483
rect 25547 25480 25559 25483
rect 26142 25480 26148 25492
rect 25547 25452 26148 25480
rect 25547 25449 25559 25452
rect 25501 25443 25559 25449
rect 26142 25440 26148 25452
rect 26200 25440 26206 25492
rect 28350 25480 28356 25492
rect 27080 25452 28356 25480
rect 21459 25384 23704 25412
rect 17368 25372 17374 25384
rect 24486 25372 24492 25424
rect 24544 25412 24550 25424
rect 24765 25415 24823 25421
rect 24765 25412 24777 25415
rect 24544 25384 24777 25412
rect 24544 25372 24550 25384
rect 24765 25381 24777 25384
rect 24811 25381 24823 25415
rect 24765 25375 24823 25381
rect 24854 25372 24860 25424
rect 24912 25412 24918 25424
rect 27080 25412 27108 25452
rect 28350 25440 28356 25452
rect 28408 25480 28414 25492
rect 28810 25480 28816 25492
rect 28408 25452 28816 25480
rect 28408 25440 28414 25452
rect 28810 25440 28816 25452
rect 28868 25440 28874 25492
rect 30926 25440 30932 25492
rect 30984 25480 30990 25492
rect 47118 25480 47124 25492
rect 30984 25452 47124 25480
rect 30984 25440 30990 25452
rect 47118 25440 47124 25452
rect 47176 25440 47182 25492
rect 24912 25384 27108 25412
rect 24912 25372 24918 25384
rect 27154 25372 27160 25424
rect 27212 25412 27218 25424
rect 38470 25412 38476 25424
rect 27212 25384 38476 25412
rect 27212 25372 27218 25384
rect 38470 25372 38476 25384
rect 38528 25372 38534 25424
rect 48041 25415 48099 25421
rect 48041 25412 48053 25415
rect 45526 25384 48053 25412
rect 13265 25347 13323 25353
rect 13265 25313 13277 25347
rect 13311 25313 13323 25347
rect 13265 25307 13323 25313
rect 13446 25304 13452 25356
rect 13504 25344 13510 25356
rect 13504 25316 14596 25344
rect 13504 25304 13510 25316
rect 11977 25279 12035 25285
rect 10928 25248 10973 25276
rect 10928 25236 10934 25248
rect 11977 25245 11989 25279
rect 12023 25245 12035 25279
rect 12250 25276 12256 25288
rect 12211 25248 12256 25276
rect 11977 25239 12035 25245
rect 12250 25236 12256 25248
rect 12308 25236 12314 25288
rect 13173 25279 13231 25285
rect 13173 25245 13185 25279
rect 13219 25276 13231 25279
rect 13906 25276 13912 25288
rect 13219 25248 13912 25276
rect 13219 25245 13231 25248
rect 13173 25239 13231 25245
rect 13906 25236 13912 25248
rect 13964 25236 13970 25288
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25276 14151 25279
rect 14182 25276 14188 25288
rect 14139 25248 14188 25276
rect 14139 25245 14151 25248
rect 14093 25239 14151 25245
rect 14182 25236 14188 25248
rect 14240 25236 14246 25288
rect 14458 25276 14464 25288
rect 14419 25248 14464 25276
rect 14458 25236 14464 25248
rect 14516 25236 14522 25288
rect 14568 25285 14596 25316
rect 15378 25304 15384 25356
rect 15436 25344 15442 25356
rect 16206 25344 16212 25356
rect 15436 25316 16212 25344
rect 15436 25304 15442 25316
rect 16206 25304 16212 25316
rect 16264 25304 16270 25356
rect 18892 25316 19380 25344
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 16476 25279 16534 25285
rect 16476 25245 16488 25279
rect 16522 25276 16534 25279
rect 16758 25276 16764 25288
rect 16522 25248 16764 25276
rect 16522 25245 16534 25248
rect 16476 25239 16534 25245
rect 16758 25236 16764 25248
rect 16816 25236 16822 25288
rect 17034 25236 17040 25288
rect 17092 25276 17098 25288
rect 18892 25276 18920 25316
rect 17092 25248 18920 25276
rect 17092 25236 17098 25248
rect 19150 25236 19156 25288
rect 19208 25276 19214 25288
rect 19245 25279 19303 25285
rect 19245 25276 19257 25279
rect 19208 25248 19257 25276
rect 19208 25236 19214 25248
rect 19245 25245 19257 25248
rect 19291 25245 19303 25279
rect 19352 25276 19380 25316
rect 19426 25304 19432 25356
rect 19484 25344 19490 25356
rect 20070 25344 20076 25356
rect 19484 25316 20076 25344
rect 19484 25304 19490 25316
rect 20070 25304 20076 25316
rect 20128 25344 20134 25356
rect 20533 25347 20591 25353
rect 20533 25344 20545 25347
rect 20128 25316 20545 25344
rect 20128 25304 20134 25316
rect 20533 25313 20545 25316
rect 20579 25313 20591 25347
rect 20533 25307 20591 25313
rect 21542 25304 21548 25356
rect 21600 25344 21606 25356
rect 23201 25347 23259 25353
rect 23201 25344 23213 25347
rect 21600 25316 23213 25344
rect 21600 25304 21606 25316
rect 23201 25313 23213 25316
rect 23247 25313 23259 25347
rect 23201 25307 23259 25313
rect 23308 25316 31754 25344
rect 19518 25276 19524 25288
rect 19352 25248 19524 25276
rect 19245 25239 19303 25245
rect 19518 25236 19524 25248
rect 19576 25236 19582 25288
rect 23308 25276 23336 25316
rect 20732 25248 23336 25276
rect 23385 25279 23443 25285
rect 20732 25208 20760 25248
rect 23385 25245 23397 25279
rect 23431 25245 23443 25279
rect 24578 25276 24584 25288
rect 24539 25248 24584 25276
rect 23385 25239 23443 25245
rect 20806 25217 20812 25220
rect 9907 25180 10640 25208
rect 13372 25180 20760 25208
rect 9907 25177 9919 25180
rect 9861 25171 9919 25177
rect 2038 25100 2044 25152
rect 2096 25140 2102 25152
rect 9122 25140 9128 25152
rect 2096 25112 9128 25140
rect 2096 25100 2102 25112
rect 9122 25100 9128 25112
rect 9180 25100 9186 25152
rect 9306 25100 9312 25152
rect 9364 25140 9370 25152
rect 13372 25140 13400 25180
rect 20800 25171 20812 25217
rect 20864 25208 20870 25220
rect 20864 25180 20900 25208
rect 21008 25180 22048 25208
rect 20806 25168 20812 25171
rect 20864 25168 20870 25180
rect 13538 25140 13544 25152
rect 9364 25112 13400 25140
rect 13499 25112 13544 25140
rect 9364 25100 9370 25112
rect 13538 25100 13544 25112
rect 13596 25100 13602 25152
rect 14366 25140 14372 25152
rect 14327 25112 14372 25140
rect 14366 25100 14372 25112
rect 14424 25100 14430 25152
rect 16574 25100 16580 25152
rect 16632 25140 16638 25152
rect 17589 25143 17647 25149
rect 17589 25140 17601 25143
rect 16632 25112 17601 25140
rect 16632 25100 16638 25112
rect 17589 25109 17601 25112
rect 17635 25109 17647 25143
rect 17589 25103 17647 25109
rect 19150 25100 19156 25152
rect 19208 25140 19214 25152
rect 19334 25140 19340 25152
rect 19208 25112 19340 25140
rect 19208 25100 19214 25112
rect 19334 25100 19340 25112
rect 19392 25100 19398 25152
rect 19978 25100 19984 25152
rect 20036 25140 20042 25152
rect 21008 25140 21036 25180
rect 20036 25112 21036 25140
rect 20036 25100 20042 25112
rect 21542 25100 21548 25152
rect 21600 25140 21606 25152
rect 21913 25143 21971 25149
rect 21913 25140 21925 25143
rect 21600 25112 21925 25140
rect 21600 25100 21606 25112
rect 21913 25109 21925 25112
rect 21959 25109 21971 25143
rect 22020 25140 22048 25180
rect 22186 25168 22192 25220
rect 22244 25208 22250 25220
rect 23109 25211 23167 25217
rect 23109 25208 23121 25211
rect 22244 25180 23121 25208
rect 22244 25168 22250 25180
rect 23109 25177 23121 25180
rect 23155 25177 23167 25211
rect 23109 25171 23167 25177
rect 23198 25168 23204 25220
rect 23256 25208 23262 25220
rect 23400 25208 23428 25239
rect 24578 25236 24584 25248
rect 24636 25236 24642 25288
rect 25317 25279 25375 25285
rect 25317 25245 25329 25279
rect 25363 25245 25375 25279
rect 26142 25276 26148 25288
rect 26103 25248 26148 25276
rect 25317 25239 25375 25245
rect 23256 25180 23428 25208
rect 25332 25208 25360 25239
rect 26142 25236 26148 25248
rect 26200 25236 26206 25288
rect 27982 25276 27988 25288
rect 27943 25248 27988 25276
rect 27982 25236 27988 25248
rect 28040 25276 28046 25288
rect 29638 25276 29644 25288
rect 28040 25248 29644 25276
rect 28040 25236 28046 25248
rect 29638 25236 29644 25248
rect 29696 25276 29702 25288
rect 29917 25279 29975 25285
rect 29917 25276 29929 25279
rect 29696 25248 29929 25276
rect 29696 25236 29702 25248
rect 29917 25245 29929 25248
rect 29963 25245 29975 25279
rect 29917 25239 29975 25245
rect 26234 25208 26240 25220
rect 25332 25180 26240 25208
rect 23256 25168 23262 25180
rect 26234 25168 26240 25180
rect 26292 25168 26298 25220
rect 27249 25211 27307 25217
rect 27249 25177 27261 25211
rect 27295 25208 27307 25211
rect 27430 25208 27436 25220
rect 27295 25180 27436 25208
rect 27295 25177 27307 25180
rect 27249 25171 27307 25177
rect 27430 25168 27436 25180
rect 27488 25208 27494 25220
rect 28258 25208 28264 25220
rect 27488 25180 28264 25208
rect 27488 25168 27494 25180
rect 28258 25168 28264 25180
rect 28316 25168 28322 25220
rect 28810 25208 28816 25220
rect 28771 25180 28816 25208
rect 28810 25168 28816 25180
rect 28868 25168 28874 25220
rect 28902 25168 28908 25220
rect 28960 25208 28966 25220
rect 31726 25208 31754 25316
rect 33502 25304 33508 25356
rect 33560 25344 33566 25356
rect 45526 25344 45554 25384
rect 48041 25381 48053 25384
rect 48087 25381 48099 25415
rect 48041 25375 48099 25381
rect 33560 25316 45554 25344
rect 33560 25304 33566 25316
rect 32309 25279 32367 25285
rect 32309 25245 32321 25279
rect 32355 25276 32367 25279
rect 32490 25276 32496 25288
rect 32355 25248 32496 25276
rect 32355 25245 32367 25248
rect 32309 25239 32367 25245
rect 32490 25236 32496 25248
rect 32548 25276 32554 25288
rect 33597 25279 33655 25285
rect 33597 25276 33609 25279
rect 32548 25248 33609 25276
rect 32548 25236 32554 25248
rect 33597 25245 33609 25248
rect 33643 25245 33655 25279
rect 33597 25239 33655 25245
rect 33686 25236 33692 25288
rect 33744 25276 33750 25288
rect 34701 25279 34759 25285
rect 34701 25276 34713 25279
rect 33744 25248 34713 25276
rect 33744 25236 33750 25248
rect 34701 25245 34713 25248
rect 34747 25245 34759 25279
rect 47854 25276 47860 25288
rect 47815 25248 47860 25276
rect 34701 25239 34759 25245
rect 47854 25236 47860 25248
rect 47912 25236 47918 25288
rect 32953 25211 33011 25217
rect 32953 25208 32965 25211
rect 28960 25180 31340 25208
rect 31726 25180 32965 25208
rect 28960 25168 28966 25180
rect 26970 25140 26976 25152
rect 22020 25112 26976 25140
rect 21913 25103 21971 25109
rect 26970 25100 26976 25112
rect 27028 25100 27034 25152
rect 30926 25100 30932 25152
rect 30984 25140 30990 25152
rect 31205 25143 31263 25149
rect 31205 25140 31217 25143
rect 30984 25112 31217 25140
rect 30984 25100 30990 25112
rect 31205 25109 31217 25112
rect 31251 25109 31263 25143
rect 31312 25140 31340 25180
rect 32953 25177 32965 25180
rect 32999 25208 33011 25211
rect 40126 25208 40132 25220
rect 32999 25180 40132 25208
rect 32999 25177 33011 25180
rect 32953 25171 33011 25177
rect 40126 25168 40132 25180
rect 40184 25168 40190 25220
rect 33502 25140 33508 25152
rect 31312 25112 33508 25140
rect 31205 25103 31263 25109
rect 33502 25100 33508 25112
rect 33560 25100 33566 25152
rect 33686 25100 33692 25152
rect 33744 25140 33750 25152
rect 33781 25143 33839 25149
rect 33781 25140 33793 25143
rect 33744 25112 33793 25140
rect 33744 25100 33750 25112
rect 33781 25109 33793 25112
rect 33827 25109 33839 25143
rect 34790 25140 34796 25152
rect 34751 25112 34796 25140
rect 33781 25103 33839 25109
rect 34790 25100 34796 25112
rect 34848 25100 34854 25152
rect 1104 25050 48852 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 48852 25050
rect 1104 24976 48852 24998
rect 9508 24908 10640 24936
rect 8849 24871 8907 24877
rect 8849 24837 8861 24871
rect 8895 24868 8907 24871
rect 9398 24868 9404 24880
rect 8895 24840 9404 24868
rect 8895 24837 8907 24840
rect 8849 24831 8907 24837
rect 9398 24828 9404 24840
rect 9456 24828 9462 24880
rect 7558 24800 7564 24812
rect 7519 24772 7564 24800
rect 7558 24760 7564 24772
rect 7616 24760 7622 24812
rect 7650 24760 7656 24812
rect 7708 24800 7714 24812
rect 7745 24803 7803 24809
rect 7745 24800 7757 24803
rect 7708 24772 7757 24800
rect 7708 24760 7714 24772
rect 7745 24769 7757 24772
rect 7791 24769 7803 24803
rect 8386 24800 8392 24812
rect 8347 24772 8392 24800
rect 7745 24763 7803 24769
rect 8386 24760 8392 24772
rect 8444 24760 8450 24812
rect 8573 24803 8631 24809
rect 8573 24769 8585 24803
rect 8619 24800 8631 24803
rect 8619 24772 8892 24800
rect 8619 24769 8631 24772
rect 8573 24763 8631 24769
rect 7929 24735 7987 24741
rect 7929 24701 7941 24735
rect 7975 24732 7987 24735
rect 8588 24732 8616 24763
rect 8754 24732 8760 24744
rect 7975 24704 8616 24732
rect 8715 24704 8760 24732
rect 7975 24701 7987 24704
rect 7929 24695 7987 24701
rect 8754 24692 8760 24704
rect 8812 24692 8818 24744
rect 8864 24732 8892 24772
rect 9214 24760 9220 24812
rect 9272 24800 9278 24812
rect 9508 24803 9536 24908
rect 9671 24809 9677 24812
rect 9565 24803 9623 24809
rect 9658 24803 9677 24809
rect 9508 24800 9577 24803
rect 9272 24775 9577 24800
rect 9272 24772 9536 24775
rect 9272 24760 9278 24772
rect 9565 24769 9577 24775
rect 9611 24772 9628 24803
rect 9611 24769 9623 24772
rect 9565 24763 9623 24769
rect 9658 24769 9670 24803
rect 9658 24763 9677 24769
rect 9671 24760 9677 24763
rect 9729 24760 9735 24812
rect 9769 24806 9827 24812
rect 9769 24772 9781 24806
rect 9815 24800 9827 24806
rect 9815 24772 9904 24800
rect 9769 24766 9827 24772
rect 8864 24724 9717 24732
rect 9876 24724 9904 24772
rect 9950 24760 9956 24812
rect 10008 24800 10014 24812
rect 10612 24809 10640 24908
rect 11974 24896 11980 24948
rect 12032 24936 12038 24948
rect 23474 24936 23480 24948
rect 12032 24908 22094 24936
rect 23435 24908 23480 24936
rect 12032 24896 12038 24908
rect 10962 24828 10968 24880
rect 11020 24868 11026 24880
rect 19978 24868 19984 24880
rect 11020 24840 19984 24868
rect 11020 24828 11026 24840
rect 19978 24828 19984 24840
rect 20036 24828 20042 24880
rect 22066 24868 22094 24908
rect 23474 24896 23480 24908
rect 23532 24896 23538 24948
rect 23584 24908 26924 24936
rect 23584 24868 23612 24908
rect 22066 24840 23612 24868
rect 23937 24871 23995 24877
rect 23937 24837 23949 24871
rect 23983 24868 23995 24871
rect 24026 24868 24032 24880
rect 23983 24840 24032 24868
rect 23983 24837 23995 24840
rect 23937 24831 23995 24837
rect 24026 24828 24032 24840
rect 24084 24828 24090 24880
rect 24121 24871 24179 24877
rect 24121 24837 24133 24871
rect 24167 24837 24179 24871
rect 26896 24868 26924 24908
rect 26970 24896 26976 24948
rect 27028 24936 27034 24948
rect 48038 24936 48044 24948
rect 27028 24908 48044 24936
rect 27028 24896 27034 24908
rect 48038 24896 48044 24908
rect 48096 24896 48102 24948
rect 32030 24868 32036 24880
rect 26896 24840 32036 24868
rect 24121 24831 24179 24837
rect 20790 24812 20848 24815
rect 10597 24803 10655 24809
rect 10008 24772 10053 24800
rect 10008 24760 10014 24772
rect 10597 24769 10609 24803
rect 10643 24800 10655 24803
rect 10643 24772 13124 24800
rect 10643 24769 10655 24772
rect 10597 24763 10655 24769
rect 8864 24704 9904 24724
rect 9689 24696 9904 24704
rect 10318 24692 10324 24744
rect 10376 24732 10382 24744
rect 10505 24735 10563 24741
rect 10505 24732 10517 24735
rect 10376 24704 10517 24732
rect 10376 24692 10382 24704
rect 10505 24701 10517 24704
rect 10551 24701 10563 24735
rect 10505 24695 10563 24701
rect 10965 24735 11023 24741
rect 10965 24701 10977 24735
rect 11011 24732 11023 24735
rect 11606 24732 11612 24744
rect 11011 24704 11612 24732
rect 11011 24701 11023 24704
rect 10965 24695 11023 24701
rect 11606 24692 11612 24704
rect 11664 24692 11670 24744
rect 13096 24732 13124 24772
rect 13170 24760 13176 24812
rect 13228 24800 13234 24812
rect 13449 24803 13507 24809
rect 13449 24800 13461 24803
rect 13228 24772 13461 24800
rect 13228 24760 13234 24772
rect 13449 24769 13461 24772
rect 13495 24769 13507 24803
rect 16574 24800 16580 24812
rect 13449 24763 13507 24769
rect 13648 24772 16580 24800
rect 13648 24732 13676 24772
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 18874 24760 18880 24812
rect 18932 24800 18938 24812
rect 18969 24803 19027 24809
rect 18969 24800 18981 24803
rect 18932 24772 18981 24800
rect 18932 24760 18938 24772
rect 18969 24769 18981 24772
rect 19015 24769 19027 24803
rect 19150 24800 19156 24812
rect 19111 24772 19156 24800
rect 18969 24763 19027 24769
rect 19150 24760 19156 24772
rect 19208 24760 19214 24812
rect 19334 24760 19340 24812
rect 19392 24800 19398 24812
rect 19392 24772 19437 24800
rect 19392 24760 19398 24772
rect 19886 24760 19892 24812
rect 19944 24800 19950 24812
rect 20790 24809 20803 24812
rect 20671 24803 20729 24809
rect 20671 24800 20683 24803
rect 19944 24772 20683 24800
rect 19944 24760 19950 24772
rect 20671 24769 20683 24772
rect 20717 24769 20729 24803
rect 20790 24775 20802 24809
rect 20790 24769 20803 24775
rect 20671 24763 20729 24769
rect 20797 24760 20803 24769
rect 20855 24760 20861 24812
rect 20901 24806 20959 24809
rect 20901 24803 21036 24806
rect 20901 24769 20913 24803
rect 20947 24778 21036 24803
rect 20947 24769 20959 24778
rect 20901 24763 20959 24769
rect 21008 24744 21036 24778
rect 21085 24803 21143 24809
rect 21085 24769 21097 24803
rect 21131 24800 21143 24803
rect 21174 24800 21180 24812
rect 21131 24772 21180 24800
rect 21131 24769 21143 24772
rect 21085 24763 21143 24769
rect 21174 24760 21180 24772
rect 21232 24760 21238 24812
rect 21358 24760 21364 24812
rect 21416 24800 21422 24812
rect 23006 24803 23064 24809
rect 23006 24800 23018 24803
rect 21416 24772 23018 24800
rect 21416 24760 21422 24772
rect 23006 24769 23018 24772
rect 23052 24769 23064 24803
rect 23293 24803 23351 24809
rect 23293 24800 23305 24803
rect 23006 24763 23064 24769
rect 23124 24772 23305 24800
rect 13096 24704 13676 24732
rect 13725 24735 13783 24741
rect 13725 24701 13737 24735
rect 13771 24732 13783 24735
rect 14366 24732 14372 24744
rect 13771 24704 14372 24732
rect 13771 24701 13783 24704
rect 13725 24695 13783 24701
rect 14366 24692 14372 24704
rect 14424 24692 14430 24744
rect 20070 24732 20076 24744
rect 17236 24704 20076 24732
rect 17236 24664 17264 24704
rect 20070 24692 20076 24704
rect 20128 24692 20134 24744
rect 20990 24692 20996 24744
rect 21048 24692 21054 24744
rect 22741 24735 22799 24741
rect 22741 24701 22753 24735
rect 22787 24732 22799 24735
rect 23124 24732 23152 24772
rect 23293 24769 23305 24772
rect 23339 24769 23351 24803
rect 23293 24763 23351 24769
rect 22787 24704 23152 24732
rect 23201 24735 23259 24741
rect 22787 24701 22799 24704
rect 22741 24695 22799 24701
rect 23201 24701 23213 24735
rect 23247 24701 23259 24735
rect 23201 24695 23259 24701
rect 20346 24664 20352 24676
rect 2746 24636 17264 24664
rect 17328 24636 20352 24664
rect 2222 24556 2228 24608
rect 2280 24596 2286 24608
rect 2746 24596 2774 24636
rect 8662 24596 8668 24608
rect 2280 24568 2774 24596
rect 8623 24568 8668 24596
rect 2280 24556 2286 24568
rect 8662 24556 8668 24568
rect 8720 24596 8726 24608
rect 9214 24596 9220 24608
rect 8720 24568 9220 24596
rect 8720 24556 8726 24568
rect 9214 24556 9220 24568
rect 9272 24556 9278 24608
rect 9309 24599 9367 24605
rect 9309 24565 9321 24599
rect 9355 24596 9367 24599
rect 10870 24596 10876 24608
rect 9355 24568 10876 24596
rect 9355 24565 9367 24568
rect 9309 24559 9367 24565
rect 10870 24556 10876 24568
rect 10928 24556 10934 24608
rect 13446 24556 13452 24608
rect 13504 24596 13510 24608
rect 13541 24599 13599 24605
rect 13541 24596 13553 24599
rect 13504 24568 13553 24596
rect 13504 24556 13510 24568
rect 13541 24565 13553 24568
rect 13587 24565 13599 24599
rect 13541 24559 13599 24565
rect 13633 24599 13691 24605
rect 13633 24565 13645 24599
rect 13679 24596 13691 24599
rect 14274 24596 14280 24608
rect 13679 24568 14280 24596
rect 13679 24565 13691 24568
rect 13633 24559 13691 24565
rect 14274 24556 14280 24568
rect 14332 24556 14338 24608
rect 15102 24556 15108 24608
rect 15160 24596 15166 24608
rect 17328 24596 17356 24636
rect 20346 24624 20352 24636
rect 20404 24624 20410 24676
rect 20441 24667 20499 24673
rect 20441 24633 20453 24667
rect 20487 24664 20499 24667
rect 20622 24664 20628 24676
rect 20487 24636 20628 24664
rect 20487 24633 20499 24636
rect 20441 24627 20499 24633
rect 20622 24624 20628 24636
rect 20680 24624 20686 24676
rect 21634 24624 21640 24676
rect 21692 24664 21698 24676
rect 21692 24636 23060 24664
rect 21692 24624 21698 24636
rect 15160 24568 17356 24596
rect 15160 24556 15166 24568
rect 18874 24556 18880 24608
rect 18932 24596 18938 24608
rect 22922 24596 22928 24608
rect 18932 24568 22928 24596
rect 18932 24556 18938 24568
rect 22922 24556 22928 24568
rect 22980 24556 22986 24608
rect 23032 24605 23060 24636
rect 23216 24608 23244 24695
rect 23308 24664 23336 24763
rect 23750 24760 23756 24812
rect 23808 24800 23814 24812
rect 24136 24800 24164 24831
rect 32030 24828 32036 24840
rect 32088 24828 32094 24880
rect 32217 24871 32275 24877
rect 32217 24837 32229 24871
rect 32263 24868 32275 24871
rect 33042 24868 33048 24880
rect 32263 24840 33048 24868
rect 32263 24837 32275 24840
rect 32217 24831 32275 24837
rect 33042 24828 33048 24840
rect 33100 24828 33106 24880
rect 23808 24772 24164 24800
rect 24949 24803 25007 24809
rect 23808 24760 23814 24772
rect 24949 24769 24961 24803
rect 24995 24769 25007 24803
rect 25682 24800 25688 24812
rect 25643 24772 25688 24800
rect 24949 24763 25007 24769
rect 24118 24692 24124 24744
rect 24176 24732 24182 24744
rect 24964 24732 24992 24763
rect 25682 24760 25688 24772
rect 25740 24760 25746 24812
rect 25866 24800 25872 24812
rect 25827 24772 25872 24800
rect 25866 24760 25872 24772
rect 25924 24760 25930 24812
rect 27065 24803 27123 24809
rect 27065 24769 27077 24803
rect 27111 24800 27123 24803
rect 27338 24800 27344 24812
rect 27111 24772 27344 24800
rect 27111 24769 27123 24772
rect 27065 24763 27123 24769
rect 27080 24732 27108 24763
rect 27338 24760 27344 24772
rect 27396 24760 27402 24812
rect 27982 24760 27988 24812
rect 28040 24800 28046 24812
rect 28077 24803 28135 24809
rect 28077 24800 28089 24803
rect 28040 24772 28089 24800
rect 28040 24760 28046 24772
rect 28077 24769 28089 24772
rect 28123 24800 28135 24803
rect 28905 24803 28963 24809
rect 28905 24800 28917 24803
rect 28123 24772 28917 24800
rect 28123 24769 28135 24772
rect 28077 24763 28135 24769
rect 28905 24769 28917 24772
rect 28951 24769 28963 24803
rect 28905 24763 28963 24769
rect 30745 24803 30803 24809
rect 30745 24769 30757 24803
rect 30791 24800 30803 24803
rect 31938 24800 31944 24812
rect 30791 24772 31944 24800
rect 30791 24769 30803 24772
rect 30745 24763 30803 24769
rect 31938 24760 31944 24772
rect 31996 24760 32002 24812
rect 32125 24803 32183 24809
rect 32125 24769 32137 24803
rect 32171 24800 32183 24803
rect 32490 24800 32496 24812
rect 32171 24772 32496 24800
rect 32171 24769 32183 24772
rect 32125 24763 32183 24769
rect 32490 24760 32496 24772
rect 32548 24760 32554 24812
rect 38010 24800 38016 24812
rect 37971 24772 38016 24800
rect 38010 24760 38016 24772
rect 38068 24760 38074 24812
rect 38286 24800 38292 24812
rect 38247 24772 38292 24800
rect 38286 24760 38292 24772
rect 38344 24760 38350 24812
rect 45646 24760 45652 24812
rect 45704 24800 45710 24812
rect 47210 24800 47216 24812
rect 45704 24772 47216 24800
rect 45704 24760 45710 24772
rect 47210 24760 47216 24772
rect 47268 24800 47274 24812
rect 47581 24803 47639 24809
rect 47581 24800 47593 24803
rect 47268 24772 47593 24800
rect 47268 24760 47274 24772
rect 47581 24769 47593 24772
rect 47627 24769 47639 24803
rect 47581 24763 47639 24769
rect 24176 24704 24348 24732
rect 24964 24704 27108 24732
rect 24176 24692 24182 24704
rect 24320 24673 24348 24704
rect 27154 24692 27160 24744
rect 27212 24732 27218 24744
rect 29273 24735 29331 24741
rect 29273 24732 29285 24735
rect 27212 24704 29285 24732
rect 27212 24692 27218 24704
rect 29273 24701 29285 24704
rect 29319 24701 29331 24735
rect 29273 24695 29331 24701
rect 29546 24692 29552 24744
rect 29604 24732 29610 24744
rect 30929 24735 30987 24741
rect 30929 24732 30941 24735
rect 29604 24704 30941 24732
rect 29604 24692 29610 24704
rect 30929 24701 30941 24704
rect 30975 24732 30987 24735
rect 31386 24732 31392 24744
rect 30975 24704 31392 24732
rect 30975 24701 30987 24704
rect 30929 24695 30987 24701
rect 31386 24692 31392 24704
rect 31444 24692 31450 24744
rect 32582 24692 32588 24744
rect 32640 24732 32646 24744
rect 32769 24735 32827 24741
rect 32769 24732 32781 24735
rect 32640 24704 32781 24732
rect 32640 24692 32646 24704
rect 32769 24701 32781 24704
rect 32815 24701 32827 24735
rect 32950 24732 32956 24744
rect 32911 24704 32956 24732
rect 32769 24695 32827 24701
rect 32950 24692 32956 24704
rect 33008 24692 33014 24744
rect 34422 24732 34428 24744
rect 34383 24704 34428 24732
rect 34422 24692 34428 24704
rect 34480 24692 34486 24744
rect 38102 24732 38108 24744
rect 38063 24704 38108 24732
rect 38102 24692 38108 24704
rect 38160 24692 38166 24744
rect 40034 24732 40040 24744
rect 39995 24704 40040 24732
rect 40034 24692 40040 24704
rect 40092 24692 40098 24744
rect 40218 24732 40224 24744
rect 40179 24704 40224 24732
rect 40218 24692 40224 24704
rect 40276 24692 40282 24744
rect 41230 24732 41236 24744
rect 41191 24704 41236 24732
rect 41230 24692 41236 24704
rect 41288 24692 41294 24744
rect 24305 24667 24363 24673
rect 23308 24636 24256 24664
rect 23017 24599 23075 24605
rect 23017 24565 23029 24599
rect 23063 24565 23075 24599
rect 23017 24559 23075 24565
rect 23198 24556 23204 24608
rect 23256 24556 23262 24608
rect 23382 24556 23388 24608
rect 23440 24596 23446 24608
rect 23658 24596 23664 24608
rect 23440 24568 23664 24596
rect 23440 24556 23446 24568
rect 23658 24556 23664 24568
rect 23716 24596 23722 24608
rect 24121 24599 24179 24605
rect 24121 24596 24133 24599
rect 23716 24568 24133 24596
rect 23716 24556 23722 24568
rect 24121 24565 24133 24568
rect 24167 24565 24179 24599
rect 24228 24596 24256 24636
rect 24305 24633 24317 24667
rect 24351 24633 24363 24667
rect 24305 24627 24363 24633
rect 24412 24636 38608 24664
rect 24412 24596 24440 24636
rect 24228 24568 24440 24596
rect 24121 24559 24179 24565
rect 24762 24556 24768 24608
rect 24820 24596 24826 24608
rect 25041 24599 25099 24605
rect 25041 24596 25053 24599
rect 24820 24568 25053 24596
rect 24820 24556 24826 24568
rect 25041 24565 25053 24568
rect 25087 24565 25099 24599
rect 25041 24559 25099 24565
rect 25866 24556 25872 24608
rect 25924 24596 25930 24608
rect 25961 24599 26019 24605
rect 25961 24596 25973 24599
rect 25924 24568 25973 24596
rect 25924 24556 25930 24568
rect 25961 24565 25973 24568
rect 26007 24565 26019 24599
rect 25961 24559 26019 24565
rect 26418 24556 26424 24608
rect 26476 24596 26482 24608
rect 27157 24599 27215 24605
rect 27157 24596 27169 24599
rect 26476 24568 27169 24596
rect 26476 24556 26482 24568
rect 27157 24565 27169 24568
rect 27203 24565 27215 24599
rect 27157 24559 27215 24565
rect 27982 24556 27988 24608
rect 28040 24596 28046 24608
rect 28169 24599 28227 24605
rect 28169 24596 28181 24599
rect 28040 24568 28181 24596
rect 28040 24556 28046 24568
rect 28169 24565 28181 24568
rect 28215 24565 28227 24599
rect 28169 24559 28227 24565
rect 29730 24556 29736 24608
rect 29788 24596 29794 24608
rect 35618 24596 35624 24608
rect 29788 24568 35624 24596
rect 29788 24556 29794 24568
rect 35618 24556 35624 24568
rect 35676 24556 35682 24608
rect 38102 24596 38108 24608
rect 38063 24568 38108 24596
rect 38102 24556 38108 24568
rect 38160 24556 38166 24608
rect 38470 24596 38476 24608
rect 38431 24568 38476 24596
rect 38470 24556 38476 24568
rect 38528 24556 38534 24608
rect 38580 24596 38608 24636
rect 38654 24624 38660 24676
rect 38712 24664 38718 24676
rect 48130 24664 48136 24676
rect 38712 24636 48136 24664
rect 38712 24624 38718 24636
rect 48130 24624 48136 24636
rect 48188 24624 48194 24676
rect 44910 24596 44916 24608
rect 38580 24568 44916 24596
rect 44910 24556 44916 24568
rect 44968 24556 44974 24608
rect 46290 24556 46296 24608
rect 46348 24596 46354 24608
rect 47029 24599 47087 24605
rect 47029 24596 47041 24599
rect 46348 24568 47041 24596
rect 46348 24556 46354 24568
rect 47029 24565 47041 24568
rect 47075 24565 47087 24599
rect 47670 24596 47676 24608
rect 47631 24568 47676 24596
rect 47029 24559 47087 24565
rect 47670 24556 47676 24568
rect 47728 24556 47734 24608
rect 1104 24506 48852 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 48852 24506
rect 1104 24432 48852 24454
rect 8386 24352 8392 24404
rect 8444 24392 8450 24404
rect 9125 24395 9183 24401
rect 9125 24392 9137 24395
rect 8444 24364 9137 24392
rect 8444 24352 8450 24364
rect 9125 24361 9137 24364
rect 9171 24392 9183 24395
rect 9950 24392 9956 24404
rect 9171 24364 9956 24392
rect 9171 24361 9183 24364
rect 9125 24355 9183 24361
rect 9950 24352 9956 24364
rect 10008 24352 10014 24404
rect 10410 24352 10416 24404
rect 10468 24392 10474 24404
rect 12894 24392 12900 24404
rect 10468 24364 12900 24392
rect 10468 24352 10474 24364
rect 12894 24352 12900 24364
rect 12952 24352 12958 24404
rect 22738 24392 22744 24404
rect 19536 24364 22744 24392
rect 7558 24284 7564 24336
rect 7616 24324 7622 24336
rect 7616 24296 12434 24324
rect 7616 24284 7622 24296
rect 9048 24200 9076 24296
rect 9582 24216 9588 24268
rect 9640 24256 9646 24268
rect 9953 24259 10011 24265
rect 9953 24256 9965 24259
rect 9640 24228 9965 24256
rect 9640 24216 9646 24228
rect 9953 24225 9965 24228
rect 9999 24256 10011 24259
rect 10318 24256 10324 24268
rect 9999 24228 10324 24256
rect 9999 24225 10011 24228
rect 9953 24219 10011 24225
rect 10318 24216 10324 24228
rect 10376 24216 10382 24268
rect 12406 24256 12434 24296
rect 19426 24256 19432 24268
rect 12406 24228 19432 24256
rect 19426 24216 19432 24228
rect 19484 24216 19490 24268
rect 1394 24188 1400 24200
rect 1355 24160 1400 24188
rect 1394 24148 1400 24160
rect 1452 24148 1458 24200
rect 9030 24188 9036 24200
rect 8991 24160 9036 24188
rect 9030 24148 9036 24160
rect 9088 24148 9094 24200
rect 9217 24191 9275 24197
rect 9217 24157 9229 24191
rect 9263 24157 9275 24191
rect 9674 24188 9680 24200
rect 9635 24160 9680 24188
rect 9217 24151 9275 24157
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 9232 24120 9260 24151
rect 9674 24148 9680 24160
rect 9732 24148 9738 24200
rect 19536 24188 19564 24364
rect 22738 24352 22744 24364
rect 22796 24352 22802 24404
rect 22830 24352 22836 24404
rect 22888 24392 22894 24404
rect 22925 24395 22983 24401
rect 22925 24392 22937 24395
rect 22888 24364 22937 24392
rect 22888 24352 22894 24364
rect 22925 24361 22937 24364
rect 22971 24361 22983 24395
rect 22925 24355 22983 24361
rect 24302 24352 24308 24404
rect 24360 24392 24366 24404
rect 24397 24395 24455 24401
rect 24397 24392 24409 24395
rect 24360 24364 24409 24392
rect 24360 24352 24366 24364
rect 24397 24361 24409 24364
rect 24443 24361 24455 24395
rect 38654 24392 38660 24404
rect 24397 24355 24455 24361
rect 24780 24364 38660 24392
rect 23014 24284 23020 24336
rect 23072 24324 23078 24336
rect 24780 24324 24808 24364
rect 38654 24352 38660 24364
rect 38712 24352 38718 24404
rect 40218 24392 40224 24404
rect 40179 24364 40224 24392
rect 40218 24352 40224 24364
rect 40276 24352 40282 24404
rect 23072 24296 24808 24324
rect 23072 24284 23078 24296
rect 32490 24284 32496 24336
rect 32548 24324 32554 24336
rect 33686 24324 33692 24336
rect 32548 24296 33692 24324
rect 32548 24284 32554 24296
rect 33686 24284 33692 24296
rect 33744 24284 33750 24336
rect 34790 24284 34796 24336
rect 34848 24324 34854 24336
rect 34848 24296 34928 24324
rect 34848 24284 34854 24296
rect 23934 24216 23940 24268
rect 23992 24256 23998 24268
rect 24486 24256 24492 24268
rect 23992 24228 24492 24256
rect 23992 24216 23998 24228
rect 24486 24216 24492 24228
rect 24544 24216 24550 24268
rect 29086 24216 29092 24268
rect 29144 24256 29150 24268
rect 34900 24265 34928 24296
rect 35618 24284 35624 24336
rect 35676 24324 35682 24336
rect 48038 24324 48044 24336
rect 35676 24296 48044 24324
rect 35676 24284 35682 24296
rect 48038 24284 48044 24296
rect 48096 24284 48102 24336
rect 34701 24259 34759 24265
rect 34701 24256 34713 24259
rect 29144 24228 34713 24256
rect 29144 24216 29150 24228
rect 34701 24225 34713 24228
rect 34747 24225 34759 24259
rect 34701 24219 34759 24225
rect 34885 24259 34943 24265
rect 34885 24225 34897 24259
rect 34931 24225 34943 24259
rect 36538 24256 36544 24268
rect 36499 24228 36544 24256
rect 34885 24219 34943 24225
rect 36538 24216 36544 24228
rect 36596 24216 36602 24268
rect 46290 24256 46296 24268
rect 46251 24228 46296 24256
rect 46290 24216 46296 24228
rect 46348 24216 46354 24268
rect 46477 24259 46535 24265
rect 46477 24225 46489 24259
rect 46523 24256 46535 24259
rect 47670 24256 47676 24268
rect 46523 24228 47676 24256
rect 46523 24225 46535 24228
rect 46477 24219 46535 24225
rect 47670 24216 47676 24228
rect 47728 24216 47734 24268
rect 48130 24256 48136 24268
rect 48091 24228 48136 24256
rect 48130 24216 48136 24228
rect 48188 24216 48194 24268
rect 12406 24160 19564 24188
rect 19705 24191 19763 24197
rect 10042 24120 10048 24132
rect 7708 24092 10048 24120
rect 7708 24080 7714 24092
rect 10042 24080 10048 24092
rect 10100 24080 10106 24132
rect 1578 24052 1584 24064
rect 1539 24024 1584 24052
rect 1578 24012 1584 24024
rect 1636 24012 1642 24064
rect 7282 24012 7288 24064
rect 7340 24052 7346 24064
rect 12406 24052 12434 24160
rect 19705 24157 19717 24191
rect 19751 24188 19763 24191
rect 21818 24188 21824 24200
rect 19751 24160 21824 24188
rect 19751 24157 19763 24160
rect 19705 24151 19763 24157
rect 21818 24148 21824 24160
rect 21876 24148 21882 24200
rect 24394 24148 24400 24200
rect 24452 24188 24458 24200
rect 24670 24188 24676 24200
rect 24452 24160 24497 24188
rect 24631 24160 24676 24188
rect 24452 24148 24458 24160
rect 24670 24148 24676 24160
rect 24728 24148 24734 24200
rect 25777 24191 25835 24197
rect 25777 24157 25789 24191
rect 25823 24188 25835 24191
rect 27614 24188 27620 24200
rect 25823 24160 27620 24188
rect 25823 24157 25835 24160
rect 25777 24151 25835 24157
rect 27614 24148 27620 24160
rect 27672 24148 27678 24200
rect 27724 24160 28120 24188
rect 12526 24080 12532 24132
rect 12584 24120 12590 24132
rect 12713 24123 12771 24129
rect 12713 24120 12725 24123
rect 12584 24092 12725 24120
rect 12584 24080 12590 24092
rect 12713 24089 12725 24092
rect 12759 24120 12771 24123
rect 13262 24120 13268 24132
rect 12759 24092 13268 24120
rect 12759 24089 12771 24092
rect 12713 24083 12771 24089
rect 13262 24080 13268 24092
rect 13320 24080 13326 24132
rect 16393 24123 16451 24129
rect 16393 24089 16405 24123
rect 16439 24089 16451 24123
rect 16574 24120 16580 24132
rect 16535 24092 16580 24120
rect 16393 24083 16451 24089
rect 7340 24024 12434 24052
rect 7340 24012 7346 24024
rect 12802 24012 12808 24064
rect 12860 24052 12866 24064
rect 12913 24055 12971 24061
rect 12913 24052 12925 24055
rect 12860 24024 12925 24052
rect 12860 24012 12866 24024
rect 12913 24021 12925 24024
rect 12959 24021 12971 24055
rect 13078 24052 13084 24064
rect 13039 24024 13084 24052
rect 12913 24015 12971 24021
rect 13078 24012 13084 24024
rect 13136 24012 13142 24064
rect 16408 24052 16436 24083
rect 16574 24080 16580 24092
rect 16632 24080 16638 24132
rect 17954 24120 17960 24132
rect 16684 24092 17960 24120
rect 16684 24052 16712 24092
rect 17954 24080 17960 24092
rect 18012 24080 18018 24132
rect 19972 24123 20030 24129
rect 19972 24089 19984 24123
rect 20018 24120 20030 24123
rect 20346 24120 20352 24132
rect 20018 24092 20352 24120
rect 20018 24089 20030 24092
rect 19972 24083 20030 24089
rect 20346 24080 20352 24092
rect 20404 24080 20410 24132
rect 21634 24120 21640 24132
rect 21595 24092 21640 24120
rect 21634 24080 21640 24092
rect 21692 24080 21698 24132
rect 21726 24080 21732 24132
rect 21784 24120 21790 24132
rect 21784 24092 22094 24120
rect 21784 24080 21790 24092
rect 16408 24024 16712 24052
rect 16761 24055 16819 24061
rect 16761 24021 16773 24055
rect 16807 24052 16819 24055
rect 17126 24052 17132 24064
rect 16807 24024 17132 24052
rect 16807 24021 16819 24024
rect 16761 24015 16819 24021
rect 17126 24012 17132 24024
rect 17184 24012 17190 24064
rect 17218 24012 17224 24064
rect 17276 24052 17282 24064
rect 20622 24052 20628 24064
rect 17276 24024 20628 24052
rect 17276 24012 17282 24024
rect 20622 24012 20628 24024
rect 20680 24012 20686 24064
rect 20714 24012 20720 24064
rect 20772 24052 20778 24064
rect 21085 24055 21143 24061
rect 21085 24052 21097 24055
rect 20772 24024 21097 24052
rect 20772 24012 20778 24024
rect 21085 24021 21097 24024
rect 21131 24021 21143 24055
rect 22066 24052 22094 24092
rect 22738 24080 22744 24132
rect 22796 24120 22802 24132
rect 22796 24092 25820 24120
rect 22796 24080 22802 24092
rect 24857 24055 24915 24061
rect 24857 24052 24869 24055
rect 22066 24024 24869 24052
rect 21085 24015 21143 24021
rect 24857 24021 24869 24024
rect 24903 24021 24915 24055
rect 25792 24052 25820 24092
rect 25866 24080 25872 24132
rect 25924 24120 25930 24132
rect 26022 24123 26080 24129
rect 26022 24120 26034 24123
rect 25924 24092 26034 24120
rect 25924 24080 25930 24092
rect 26022 24089 26034 24092
rect 26068 24089 26080 24123
rect 27724 24120 27752 24160
rect 27890 24129 27896 24132
rect 26022 24083 26080 24089
rect 26988 24092 27752 24120
rect 26988 24052 27016 24092
rect 27884 24083 27896 24129
rect 27948 24120 27954 24132
rect 28092 24120 28120 24160
rect 28166 24148 28172 24200
rect 28224 24188 28230 24200
rect 29638 24188 29644 24200
rect 28224 24160 29500 24188
rect 29599 24160 29644 24188
rect 28224 24148 28230 24160
rect 28350 24120 28356 24132
rect 27948 24092 27984 24120
rect 28092 24092 28356 24120
rect 27890 24080 27896 24083
rect 27948 24080 27954 24092
rect 28350 24080 28356 24092
rect 28408 24080 28414 24132
rect 29472 24120 29500 24160
rect 29638 24148 29644 24160
rect 29696 24148 29702 24200
rect 30745 24191 30803 24197
rect 30745 24188 30757 24191
rect 29748 24160 30757 24188
rect 29748 24120 29776 24160
rect 30745 24157 30757 24160
rect 30791 24157 30803 24191
rect 31386 24188 31392 24200
rect 31347 24160 31392 24188
rect 30745 24151 30803 24157
rect 31386 24148 31392 24160
rect 31444 24148 31450 24200
rect 32858 24148 32864 24200
rect 32916 24188 32922 24200
rect 33229 24191 33287 24197
rect 33229 24188 33241 24191
rect 32916 24160 33241 24188
rect 32916 24148 32922 24160
rect 33229 24157 33241 24160
rect 33275 24157 33287 24191
rect 33686 24188 33692 24200
rect 33647 24160 33692 24188
rect 33229 24151 33287 24157
rect 33686 24148 33692 24160
rect 33744 24148 33750 24200
rect 40126 24188 40132 24200
rect 40087 24160 40132 24188
rect 40126 24148 40132 24160
rect 40184 24148 40190 24200
rect 30006 24120 30012 24132
rect 28644 24092 29408 24120
rect 29472 24092 29776 24120
rect 29967 24092 30012 24120
rect 27154 24052 27160 24064
rect 25792 24024 27016 24052
rect 27067 24024 27160 24052
rect 24857 24015 24915 24021
rect 27154 24012 27160 24024
rect 27212 24052 27218 24064
rect 28644 24052 28672 24092
rect 27212 24024 28672 24052
rect 27212 24012 27218 24024
rect 28994 24012 29000 24064
rect 29052 24052 29058 24064
rect 29380 24052 29408 24092
rect 30006 24080 30012 24092
rect 30064 24080 30070 24132
rect 30837 24123 30895 24129
rect 30837 24089 30849 24123
rect 30883 24120 30895 24123
rect 31573 24123 31631 24129
rect 31573 24120 31585 24123
rect 30883 24092 31585 24120
rect 30883 24089 30895 24092
rect 30837 24083 30895 24089
rect 31573 24089 31585 24092
rect 31619 24089 31631 24123
rect 40034 24120 40040 24132
rect 31573 24083 31631 24089
rect 31680 24092 40040 24120
rect 31680 24052 31708 24092
rect 40034 24080 40040 24092
rect 40092 24080 40098 24132
rect 29052 24024 29097 24052
rect 29380 24024 31708 24052
rect 29052 24012 29058 24024
rect 33410 24012 33416 24064
rect 33468 24052 33474 24064
rect 33781 24055 33839 24061
rect 33781 24052 33793 24055
rect 33468 24024 33793 24052
rect 33468 24012 33474 24024
rect 33781 24021 33793 24024
rect 33827 24021 33839 24055
rect 33781 24015 33839 24021
rect 1104 23962 48852 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 48852 23962
rect 1104 23888 48852 23910
rect 1578 23808 1584 23860
rect 1636 23848 1642 23860
rect 12618 23848 12624 23860
rect 1636 23820 12624 23848
rect 1636 23808 1642 23820
rect 12618 23808 12624 23820
rect 12676 23808 12682 23860
rect 12713 23851 12771 23857
rect 12713 23817 12725 23851
rect 12759 23848 12771 23851
rect 12894 23848 12900 23860
rect 12759 23820 12900 23848
rect 12759 23817 12771 23820
rect 12713 23811 12771 23817
rect 12894 23808 12900 23820
rect 12952 23848 12958 23860
rect 13722 23848 13728 23860
rect 12952 23820 13728 23848
rect 12952 23808 12958 23820
rect 13722 23808 13728 23820
rect 13780 23808 13786 23860
rect 18506 23848 18512 23860
rect 14108 23820 16988 23848
rect 14108 23780 14136 23820
rect 14274 23780 14280 23792
rect 2746 23752 14136 23780
rect 14235 23752 14280 23780
rect 2314 23536 2320 23588
rect 2372 23576 2378 23588
rect 2746 23576 2774 23752
rect 14274 23740 14280 23752
rect 14332 23740 14338 23792
rect 7374 23712 7380 23724
rect 7335 23684 7380 23712
rect 7374 23672 7380 23684
rect 7432 23672 7438 23724
rect 9490 23672 9496 23724
rect 9548 23712 9554 23724
rect 9677 23715 9735 23721
rect 9677 23712 9689 23715
rect 9548 23684 9689 23712
rect 9548 23672 9554 23684
rect 9677 23681 9689 23684
rect 9723 23681 9735 23715
rect 9677 23675 9735 23681
rect 9769 23715 9827 23721
rect 9769 23681 9781 23715
rect 9815 23712 9827 23715
rect 10410 23712 10416 23724
rect 9815 23684 10416 23712
rect 9815 23681 9827 23684
rect 9769 23675 9827 23681
rect 10410 23672 10416 23684
rect 10468 23672 10474 23724
rect 11698 23712 11704 23724
rect 11659 23684 11704 23712
rect 11698 23672 11704 23684
rect 11756 23672 11762 23724
rect 12526 23672 12532 23724
rect 12584 23712 12590 23724
rect 12584 23684 12629 23712
rect 12584 23672 12590 23684
rect 12802 23672 12808 23724
rect 12860 23712 12866 23724
rect 12860 23684 12905 23712
rect 12860 23672 12866 23684
rect 13354 23672 13360 23724
rect 13412 23712 13418 23724
rect 13449 23715 13507 23721
rect 13449 23712 13461 23715
rect 13412 23684 13461 23712
rect 13412 23672 13418 23684
rect 13449 23681 13461 23684
rect 13495 23681 13507 23715
rect 13449 23675 13507 23681
rect 14550 23672 14556 23724
rect 14608 23712 14614 23724
rect 16960 23721 16988 23820
rect 17512 23820 18512 23848
rect 17218 23780 17224 23792
rect 17052 23752 17224 23780
rect 17052 23721 17080 23752
rect 17218 23740 17224 23752
rect 17276 23740 17282 23792
rect 17512 23724 17540 23820
rect 18506 23808 18512 23820
rect 18564 23808 18570 23860
rect 20346 23848 20352 23860
rect 20307 23820 20352 23848
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20990 23848 20996 23860
rect 20456 23820 20996 23848
rect 17954 23740 17960 23792
rect 18012 23780 18018 23792
rect 19150 23780 19156 23792
rect 18012 23752 19156 23780
rect 18012 23740 18018 23752
rect 19150 23740 19156 23752
rect 19208 23780 19214 23792
rect 19245 23783 19303 23789
rect 19245 23780 19257 23783
rect 19208 23752 19257 23780
rect 19208 23740 19214 23752
rect 19245 23749 19257 23752
rect 19291 23749 19303 23783
rect 19426 23780 19432 23792
rect 19387 23752 19432 23780
rect 19245 23743 19303 23749
rect 19426 23740 19432 23752
rect 19484 23740 19490 23792
rect 19613 23783 19671 23789
rect 19613 23749 19625 23783
rect 19659 23780 19671 23783
rect 20456 23780 20484 23820
rect 20990 23808 20996 23820
rect 21048 23808 21054 23860
rect 23109 23851 23167 23857
rect 23109 23817 23121 23851
rect 23155 23848 23167 23851
rect 23290 23848 23296 23860
rect 23155 23820 23296 23848
rect 23155 23817 23167 23820
rect 23109 23811 23167 23817
rect 23290 23808 23296 23820
rect 23348 23808 23354 23860
rect 25777 23851 25835 23857
rect 25777 23817 25789 23851
rect 25823 23848 25835 23851
rect 25866 23848 25872 23860
rect 25823 23820 25872 23848
rect 25823 23817 25835 23820
rect 25777 23811 25835 23817
rect 25866 23808 25872 23820
rect 25924 23808 25930 23860
rect 27341 23851 27399 23857
rect 27341 23848 27353 23851
rect 26252 23820 27353 23848
rect 23014 23780 23020 23792
rect 19659 23752 20484 23780
rect 20548 23752 23020 23780
rect 19659 23749 19671 23752
rect 19613 23743 19671 23749
rect 16945 23715 17003 23721
rect 14608 23684 14653 23712
rect 14608 23672 14614 23684
rect 16945 23681 16957 23715
rect 16991 23681 17003 23715
rect 16945 23675 17003 23681
rect 17037 23715 17095 23721
rect 17037 23681 17049 23715
rect 17083 23681 17095 23715
rect 17037 23675 17095 23681
rect 17126 23672 17132 23724
rect 17184 23712 17190 23724
rect 17313 23715 17371 23721
rect 17184 23684 17229 23712
rect 17184 23672 17190 23684
rect 17313 23681 17325 23715
rect 17359 23712 17371 23715
rect 17494 23712 17500 23724
rect 17359 23684 17500 23712
rect 17359 23681 17371 23684
rect 17313 23675 17371 23681
rect 17494 23672 17500 23684
rect 17552 23672 17558 23724
rect 18046 23672 18052 23724
rect 18104 23721 18110 23724
rect 18104 23715 18153 23721
rect 18104 23681 18107 23715
rect 18141 23681 18153 23715
rect 18104 23675 18153 23681
rect 18214 23715 18272 23721
rect 18214 23681 18226 23715
rect 18260 23681 18272 23715
rect 18214 23675 18272 23681
rect 18104 23672 18110 23675
rect 7558 23644 7564 23656
rect 7519 23616 7564 23644
rect 7558 23604 7564 23616
rect 7616 23604 7622 23656
rect 9122 23644 9128 23656
rect 9083 23616 9128 23644
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9582 23604 9588 23656
rect 9640 23644 9646 23656
rect 9953 23647 10011 23653
rect 9953 23644 9965 23647
rect 9640 23616 9965 23644
rect 9640 23604 9646 23616
rect 9953 23613 9965 23616
rect 9999 23613 10011 23647
rect 11606 23644 11612 23656
rect 11567 23616 11612 23644
rect 9953 23607 10011 23613
rect 11606 23604 11612 23616
rect 11664 23604 11670 23656
rect 13538 23644 13544 23656
rect 13499 23616 13544 23644
rect 13538 23604 13544 23616
rect 13596 23604 13602 23656
rect 14369 23647 14427 23653
rect 14369 23644 14381 23647
rect 13832 23616 14381 23644
rect 11974 23576 11980 23588
rect 2372 23548 2774 23576
rect 3896 23548 11980 23576
rect 2372 23536 2378 23548
rect 2038 23508 2044 23520
rect 1999 23480 2044 23508
rect 2038 23468 2044 23480
rect 2096 23468 2102 23520
rect 2682 23468 2688 23520
rect 2740 23508 2746 23520
rect 3896 23508 3924 23548
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 12069 23579 12127 23585
rect 12069 23545 12081 23579
rect 12115 23576 12127 23579
rect 12618 23576 12624 23588
rect 12115 23548 12624 23576
rect 12115 23545 12127 23548
rect 12069 23539 12127 23545
rect 12618 23536 12624 23548
rect 12676 23536 12682 23588
rect 13832 23585 13860 23616
rect 14369 23613 14381 23616
rect 14415 23613 14427 23647
rect 14369 23607 14427 23613
rect 17218 23604 17224 23656
rect 17276 23644 17282 23656
rect 18228 23644 18256 23675
rect 18322 23672 18328 23724
rect 18380 23712 18386 23724
rect 18506 23712 18512 23724
rect 18380 23684 18425 23712
rect 18467 23684 18512 23712
rect 18380 23672 18386 23684
rect 18506 23672 18512 23684
rect 18564 23712 18570 23724
rect 20070 23712 20076 23724
rect 18564 23684 20076 23712
rect 18564 23672 18570 23684
rect 20070 23672 20076 23684
rect 20128 23672 20134 23724
rect 20548 23715 20576 23752
rect 23014 23740 23020 23752
rect 23072 23740 23078 23792
rect 20625 23715 20683 23721
rect 20548 23687 20637 23715
rect 20625 23681 20637 23687
rect 20671 23681 20683 23715
rect 20625 23675 20683 23681
rect 20714 23715 20772 23721
rect 20714 23681 20726 23715
rect 20760 23681 20772 23715
rect 20714 23675 20772 23681
rect 17276 23616 18256 23644
rect 17276 23604 17282 23616
rect 18414 23604 18420 23656
rect 18472 23644 18478 23656
rect 20346 23644 20352 23656
rect 18472 23616 20352 23644
rect 18472 23604 18478 23616
rect 20346 23604 20352 23616
rect 20404 23604 20410 23656
rect 13817 23579 13875 23585
rect 13817 23545 13829 23579
rect 13863 23545 13875 23579
rect 13817 23539 13875 23545
rect 13924 23548 16804 23576
rect 9858 23508 9864 23520
rect 2740 23480 3924 23508
rect 9819 23480 9864 23508
rect 2740 23468 2746 23480
rect 9858 23468 9864 23480
rect 9916 23468 9922 23520
rect 12526 23508 12532 23520
rect 12487 23480 12532 23508
rect 12526 23468 12532 23480
rect 12584 23468 12590 23520
rect 12710 23468 12716 23520
rect 12768 23508 12774 23520
rect 13924 23508 13952 23548
rect 14458 23508 14464 23520
rect 12768 23480 13952 23508
rect 14419 23480 14464 23508
rect 12768 23468 12774 23480
rect 14458 23468 14464 23480
rect 14516 23468 14522 23520
rect 14734 23508 14740 23520
rect 14695 23480 14740 23508
rect 14734 23468 14740 23480
rect 14792 23468 14798 23520
rect 16666 23508 16672 23520
rect 16627 23480 16672 23508
rect 16666 23468 16672 23480
rect 16724 23468 16730 23520
rect 16776 23508 16804 23548
rect 20622 23536 20628 23588
rect 20680 23576 20686 23588
rect 20732 23576 20760 23675
rect 20806 23672 20812 23724
rect 20864 23721 20870 23724
rect 20864 23712 20872 23721
rect 20993 23715 21051 23721
rect 20864 23684 20909 23712
rect 20864 23675 20872 23684
rect 20993 23681 21005 23715
rect 21039 23699 21051 23715
rect 21174 23712 21180 23724
rect 21100 23699 21180 23712
rect 21039 23684 21180 23699
rect 21039 23681 21128 23684
rect 20993 23675 21128 23681
rect 20864 23672 20870 23675
rect 21008 23671 21128 23675
rect 21174 23672 21180 23684
rect 21232 23672 21238 23724
rect 23201 23715 23259 23721
rect 23201 23681 23213 23715
rect 23247 23681 23259 23715
rect 23201 23675 23259 23681
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23712 23351 23715
rect 23339 23684 23428 23712
rect 23339 23681 23351 23684
rect 23293 23675 23351 23681
rect 23014 23604 23020 23656
rect 23072 23644 23078 23656
rect 23216 23644 23244 23675
rect 23072 23616 23244 23644
rect 23400 23644 23428 23684
rect 23842 23672 23848 23724
rect 23900 23712 23906 23724
rect 24121 23715 24179 23721
rect 24121 23712 24133 23715
rect 23900 23684 24133 23712
rect 23900 23672 23906 23684
rect 24121 23681 24133 23684
rect 24167 23681 24179 23715
rect 24121 23675 24179 23681
rect 24213 23715 24271 23721
rect 24213 23681 24225 23715
rect 24259 23681 24271 23715
rect 24213 23675 24271 23681
rect 23750 23644 23756 23656
rect 23400 23616 23756 23644
rect 23072 23604 23078 23616
rect 23750 23604 23756 23616
rect 23808 23644 23814 23656
rect 24228 23644 24256 23675
rect 24394 23672 24400 23724
rect 24452 23712 24458 23724
rect 24673 23715 24731 23721
rect 24673 23712 24685 23715
rect 24452 23684 24685 23712
rect 24452 23672 24458 23684
rect 24673 23681 24685 23684
rect 24719 23681 24731 23715
rect 24673 23675 24731 23681
rect 25866 23672 25872 23724
rect 25924 23712 25930 23724
rect 26252 23721 26280 23820
rect 27341 23817 27353 23820
rect 27387 23817 27399 23851
rect 27890 23848 27896 23860
rect 27851 23820 27896 23848
rect 27341 23811 27399 23817
rect 27890 23808 27896 23820
rect 27948 23808 27954 23860
rect 28350 23808 28356 23860
rect 28408 23848 28414 23860
rect 30006 23848 30012 23860
rect 28408 23820 30012 23848
rect 28408 23808 28414 23820
rect 30006 23808 30012 23820
rect 30064 23808 30070 23860
rect 30374 23808 30380 23860
rect 30432 23848 30438 23860
rect 31570 23848 31576 23860
rect 30432 23820 31576 23848
rect 30432 23808 30438 23820
rect 31570 23808 31576 23820
rect 31628 23808 31634 23860
rect 32677 23851 32735 23857
rect 32677 23817 32689 23851
rect 32723 23848 32735 23851
rect 32950 23848 32956 23860
rect 32723 23820 32956 23848
rect 32723 23817 32735 23820
rect 32677 23811 32735 23817
rect 32950 23808 32956 23820
rect 33008 23808 33014 23860
rect 48038 23848 48044 23860
rect 47999 23820 48044 23848
rect 48038 23808 48044 23820
rect 48096 23808 48102 23860
rect 26602 23740 26608 23792
rect 26660 23780 26666 23792
rect 47302 23780 47308 23792
rect 26660 23752 47308 23780
rect 26660 23740 26666 23752
rect 47302 23740 47308 23752
rect 47360 23740 47366 23792
rect 47946 23780 47952 23792
rect 47907 23752 47952 23780
rect 47946 23740 47952 23752
rect 48004 23740 48010 23792
rect 26007 23715 26065 23721
rect 26007 23712 26019 23715
rect 25924 23684 26019 23712
rect 25924 23672 25930 23684
rect 26007 23681 26019 23684
rect 26053 23681 26065 23715
rect 26007 23675 26065 23681
rect 26142 23715 26200 23721
rect 26142 23681 26154 23715
rect 26188 23681 26200 23715
rect 26142 23675 26200 23681
rect 26237 23715 26295 23721
rect 26237 23681 26249 23715
rect 26283 23681 26295 23715
rect 26237 23675 26295 23681
rect 26421 23715 26479 23721
rect 26421 23681 26433 23715
rect 26467 23712 26479 23715
rect 26786 23712 26792 23724
rect 26467 23684 26792 23712
rect 26467 23681 26479 23684
rect 26421 23675 26479 23681
rect 23808 23616 24256 23644
rect 24581 23647 24639 23653
rect 23808 23604 23814 23616
rect 24581 23613 24593 23647
rect 24627 23644 24639 23647
rect 24627 23616 24716 23644
rect 24627 23613 24639 23616
rect 24581 23607 24639 23613
rect 24688 23588 24716 23616
rect 25774 23604 25780 23656
rect 25832 23644 25838 23656
rect 26160 23644 26188 23675
rect 26786 23672 26792 23684
rect 26844 23672 26850 23724
rect 26970 23712 26976 23724
rect 26931 23684 26976 23712
rect 26970 23672 26976 23684
rect 27028 23672 27034 23724
rect 27154 23712 27160 23724
rect 27115 23684 27160 23712
rect 27154 23672 27160 23684
rect 27212 23672 27218 23724
rect 27798 23672 27804 23724
rect 27856 23712 27862 23724
rect 28169 23715 28227 23721
rect 28169 23712 28181 23715
rect 27856 23684 28181 23712
rect 27856 23672 27862 23684
rect 28169 23681 28181 23684
rect 28215 23681 28227 23715
rect 28169 23675 28227 23681
rect 28261 23715 28319 23721
rect 28261 23681 28273 23715
rect 28307 23681 28319 23715
rect 28261 23675 28319 23681
rect 28074 23644 28080 23656
rect 25832 23616 28080 23644
rect 25832 23604 25838 23616
rect 28074 23604 28080 23616
rect 28132 23644 28138 23656
rect 28276 23644 28304 23675
rect 28350 23672 28356 23724
rect 28408 23712 28414 23724
rect 28537 23715 28595 23721
rect 28408 23684 28453 23712
rect 28408 23672 28414 23684
rect 28537 23681 28549 23715
rect 28583 23681 28595 23715
rect 29362 23712 29368 23724
rect 29323 23684 29368 23712
rect 28537 23675 28595 23681
rect 28132 23616 28304 23644
rect 28132 23604 28138 23616
rect 21910 23576 21916 23588
rect 20680 23548 21916 23576
rect 20680 23536 20686 23548
rect 21910 23536 21916 23548
rect 21968 23536 21974 23588
rect 22922 23576 22928 23588
rect 22883 23548 22928 23576
rect 22922 23536 22928 23548
rect 22980 23536 22986 23588
rect 24670 23536 24676 23588
rect 24728 23536 24734 23588
rect 26786 23536 26792 23588
rect 26844 23576 26850 23588
rect 28552 23576 28580 23675
rect 29362 23672 29368 23684
rect 29420 23672 29426 23724
rect 29549 23715 29607 23721
rect 29549 23681 29561 23715
rect 29595 23712 29607 23715
rect 30282 23712 30288 23724
rect 29595 23684 30288 23712
rect 29595 23681 29607 23684
rect 29549 23675 29607 23681
rect 30282 23672 30288 23684
rect 30340 23672 30346 23724
rect 30466 23721 30472 23724
rect 30460 23675 30472 23721
rect 30524 23712 30530 23724
rect 30524 23684 30560 23712
rect 30466 23672 30472 23675
rect 30524 23672 30530 23684
rect 32490 23672 32496 23724
rect 32548 23712 32554 23724
rect 32585 23715 32643 23721
rect 32585 23712 32597 23715
rect 32548 23684 32597 23712
rect 32548 23672 32554 23684
rect 32585 23681 32597 23684
rect 32631 23681 32643 23715
rect 32585 23675 32643 23681
rect 30190 23644 30196 23656
rect 30151 23616 30196 23644
rect 30190 23604 30196 23616
rect 30248 23604 30254 23656
rect 33226 23644 33232 23656
rect 33187 23616 33232 23644
rect 33226 23604 33232 23616
rect 33284 23604 33290 23656
rect 33410 23644 33416 23656
rect 33371 23616 33416 23644
rect 33410 23604 33416 23616
rect 33468 23604 33474 23656
rect 33778 23644 33784 23656
rect 33739 23616 33784 23644
rect 33778 23604 33784 23616
rect 33836 23604 33842 23656
rect 28902 23576 28908 23588
rect 26844 23548 28908 23576
rect 26844 23536 26850 23548
rect 28902 23536 28908 23548
rect 28960 23536 28966 23588
rect 17678 23508 17684 23520
rect 16776 23480 17684 23508
rect 17678 23468 17684 23480
rect 17736 23468 17742 23520
rect 17862 23508 17868 23520
rect 17823 23480 17868 23508
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 19426 23468 19432 23520
rect 19484 23508 19490 23520
rect 21542 23508 21548 23520
rect 19484 23480 21548 23508
rect 19484 23468 19490 23480
rect 21542 23468 21548 23480
rect 21600 23468 21606 23520
rect 23477 23511 23535 23517
rect 23477 23477 23489 23511
rect 23523 23508 23535 23511
rect 23658 23508 23664 23520
rect 23523 23480 23664 23508
rect 23523 23477 23535 23480
rect 23477 23471 23535 23477
rect 23658 23468 23664 23480
rect 23716 23468 23722 23520
rect 26234 23468 26240 23520
rect 26292 23508 26298 23520
rect 29546 23508 29552 23520
rect 26292 23480 29552 23508
rect 26292 23468 26298 23480
rect 29546 23468 29552 23480
rect 29604 23468 29610 23520
rect 29733 23511 29791 23517
rect 29733 23477 29745 23511
rect 29779 23508 29791 23511
rect 30374 23508 30380 23520
rect 29779 23480 30380 23508
rect 29779 23477 29791 23480
rect 29733 23471 29791 23477
rect 30374 23468 30380 23480
rect 30432 23468 30438 23520
rect 1104 23418 48852 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 48852 23418
rect 1104 23344 48852 23366
rect 7558 23264 7564 23316
rect 7616 23304 7622 23316
rect 7837 23307 7895 23313
rect 7837 23304 7849 23307
rect 7616 23276 7849 23304
rect 7616 23264 7622 23276
rect 7837 23273 7849 23276
rect 7883 23273 7895 23307
rect 9490 23304 9496 23316
rect 9403 23276 9496 23304
rect 7837 23267 7895 23273
rect 9490 23264 9496 23276
rect 9548 23264 9554 23316
rect 9674 23304 9680 23316
rect 9635 23276 9680 23304
rect 9674 23264 9680 23276
rect 9732 23264 9738 23316
rect 9766 23264 9772 23316
rect 9824 23304 9830 23316
rect 10689 23307 10747 23313
rect 9824 23276 10456 23304
rect 9824 23264 9830 23276
rect 2498 23196 2504 23248
rect 2556 23236 2562 23248
rect 4706 23236 4712 23248
rect 2556 23208 4712 23236
rect 2556 23196 2562 23208
rect 4706 23196 4712 23208
rect 4764 23236 4770 23248
rect 9508 23236 9536 23264
rect 10318 23236 10324 23248
rect 4764 23208 6684 23236
rect 9508 23208 10324 23236
rect 4764 23196 4770 23208
rect 1397 23171 1455 23177
rect 1397 23137 1409 23171
rect 1443 23168 1455 23171
rect 2038 23168 2044 23180
rect 1443 23140 2044 23168
rect 1443 23137 1455 23140
rect 1397 23131 1455 23137
rect 2038 23128 2044 23140
rect 2096 23128 2102 23180
rect 2774 23128 2780 23180
rect 2832 23168 2838 23180
rect 2832 23140 2877 23168
rect 2832 23128 2838 23140
rect 1581 23035 1639 23041
rect 1581 23001 1593 23035
rect 1627 23032 1639 23035
rect 2590 23032 2596 23044
rect 1627 23004 2596 23032
rect 1627 23001 1639 23004
rect 1581 22995 1639 23001
rect 2590 22992 2596 23004
rect 2648 22992 2654 23044
rect 6656 22964 6684 23208
rect 10318 23196 10324 23208
rect 10376 23196 10382 23248
rect 10428 23236 10456 23276
rect 10689 23273 10701 23307
rect 10735 23304 10747 23307
rect 11606 23304 11612 23316
rect 10735 23276 11612 23304
rect 10735 23273 10747 23276
rect 10689 23267 10747 23273
rect 11606 23264 11612 23276
rect 11664 23264 11670 23316
rect 12526 23304 12532 23316
rect 12487 23276 12532 23304
rect 12526 23264 12532 23276
rect 12584 23264 12590 23316
rect 12986 23304 12992 23316
rect 12947 23276 12992 23304
rect 12986 23264 12992 23276
rect 13044 23264 13050 23316
rect 14274 23304 14280 23316
rect 14235 23276 14280 23304
rect 14274 23264 14280 23276
rect 14332 23264 14338 23316
rect 14458 23304 14464 23316
rect 14419 23276 14464 23304
rect 14458 23264 14464 23276
rect 14516 23264 14522 23316
rect 15580 23276 22094 23304
rect 15580 23236 15608 23276
rect 10428 23208 15608 23236
rect 16574 23196 16580 23248
rect 16632 23236 16638 23248
rect 16945 23239 17003 23245
rect 16945 23236 16957 23239
rect 16632 23208 16957 23236
rect 16632 23196 16638 23208
rect 16945 23205 16957 23208
rect 16991 23205 17003 23239
rect 16945 23199 17003 23205
rect 18049 23239 18107 23245
rect 18049 23205 18061 23239
rect 18095 23236 18107 23239
rect 18322 23236 18328 23248
rect 18095 23208 18328 23236
rect 18095 23205 18107 23208
rect 18049 23199 18107 23205
rect 18322 23196 18328 23208
rect 18380 23196 18386 23248
rect 20533 23239 20591 23245
rect 20533 23205 20545 23239
rect 20579 23236 20591 23239
rect 20806 23236 20812 23248
rect 20579 23208 20812 23236
rect 20579 23205 20591 23208
rect 20533 23199 20591 23205
rect 20806 23196 20812 23208
rect 20864 23196 20870 23248
rect 22066 23236 22094 23276
rect 23934 23264 23940 23316
rect 23992 23304 23998 23316
rect 24302 23304 24308 23316
rect 23992 23276 24308 23304
rect 23992 23264 23998 23276
rect 24302 23264 24308 23276
rect 24360 23304 24366 23316
rect 24397 23307 24455 23313
rect 24397 23304 24409 23307
rect 24360 23276 24409 23304
rect 24360 23264 24366 23276
rect 24397 23273 24409 23276
rect 24443 23273 24455 23307
rect 24397 23267 24455 23273
rect 25682 23264 25688 23316
rect 25740 23304 25746 23316
rect 25958 23304 25964 23316
rect 25740 23276 25964 23304
rect 25740 23264 25746 23276
rect 25958 23264 25964 23276
rect 26016 23264 26022 23316
rect 28350 23264 28356 23316
rect 28408 23304 28414 23316
rect 28813 23307 28871 23313
rect 28813 23304 28825 23307
rect 28408 23276 28825 23304
rect 28408 23264 28414 23276
rect 28813 23273 28825 23276
rect 28859 23273 28871 23307
rect 28813 23267 28871 23273
rect 29917 23307 29975 23313
rect 29917 23273 29929 23307
rect 29963 23304 29975 23307
rect 30466 23304 30472 23316
rect 29963 23276 30472 23304
rect 29963 23273 29975 23276
rect 29917 23267 29975 23273
rect 30466 23264 30472 23276
rect 30524 23264 30530 23316
rect 24857 23239 24915 23245
rect 22066 23208 24808 23236
rect 10410 23168 10416 23180
rect 9324 23140 10416 23168
rect 7742 23100 7748 23112
rect 7703 23072 7748 23100
rect 7742 23060 7748 23072
rect 7800 23100 7806 23112
rect 8018 23100 8024 23112
rect 7800 23072 8024 23100
rect 7800 23060 7806 23072
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 9324 23109 9352 23140
rect 10410 23128 10416 23140
rect 10468 23128 10474 23180
rect 12618 23168 12624 23180
rect 12579 23140 12624 23168
rect 12618 23128 12624 23140
rect 12676 23128 12682 23180
rect 14734 23168 14740 23180
rect 12728 23140 14740 23168
rect 9309 23103 9367 23109
rect 9309 23069 9321 23103
rect 9355 23069 9367 23103
rect 9309 23063 9367 23069
rect 9493 23103 9551 23109
rect 9493 23069 9505 23103
rect 9539 23069 9551 23103
rect 10318 23100 10324 23112
rect 10279 23072 10324 23100
rect 9493 23063 9551 23069
rect 9508 23032 9536 23063
rect 10318 23060 10324 23072
rect 10376 23060 10382 23112
rect 12529 23103 12587 23109
rect 12529 23069 12541 23103
rect 12575 23100 12587 23103
rect 12728 23100 12756 23140
rect 14734 23128 14740 23140
rect 14792 23128 14798 23180
rect 24026 23168 24032 23180
rect 22940 23140 24032 23168
rect 22940 23112 22968 23140
rect 12575 23072 12756 23100
rect 12805 23103 12863 23109
rect 12575 23069 12587 23072
rect 12529 23063 12587 23069
rect 12805 23069 12817 23103
rect 12851 23100 12863 23103
rect 13078 23100 13084 23112
rect 12851 23072 13084 23100
rect 12851 23069 12863 23072
rect 12805 23063 12863 23069
rect 13078 23060 13084 23072
rect 13136 23060 13142 23112
rect 15562 23100 15568 23112
rect 14016 23072 15424 23100
rect 15523 23072 15568 23100
rect 9582 23032 9588 23044
rect 9495 23004 9588 23032
rect 9582 22992 9588 23004
rect 9640 23032 9646 23044
rect 14016 23032 14044 23072
rect 9640 23004 14044 23032
rect 9640 22992 9646 23004
rect 14090 22992 14096 23044
rect 14148 23041 14154 23044
rect 14366 23041 14372 23044
rect 14148 23035 14177 23041
rect 14165 23001 14177 23035
rect 14309 23035 14372 23041
rect 14309 23032 14321 23035
rect 14148 22995 14177 23001
rect 14292 23001 14321 23032
rect 14355 23001 14372 23035
rect 14292 22995 14372 23001
rect 14148 22992 14154 22995
rect 9766 22964 9772 22976
rect 6656 22936 9772 22964
rect 9766 22924 9772 22936
rect 9824 22924 9830 22976
rect 13630 22924 13636 22976
rect 13688 22964 13694 22976
rect 14292 22964 14320 22995
rect 14366 22992 14372 22995
rect 14424 22992 14430 23044
rect 15396 23032 15424 23072
rect 15562 23060 15568 23072
rect 15620 23060 15626 23112
rect 15832 23103 15890 23109
rect 15832 23069 15844 23103
rect 15878 23100 15890 23103
rect 16666 23100 16672 23112
rect 15878 23072 16672 23100
rect 15878 23069 15890 23072
rect 15832 23063 15890 23069
rect 16666 23060 16672 23072
rect 16724 23060 16730 23112
rect 17865 23103 17923 23109
rect 17865 23100 17877 23103
rect 16776 23072 17877 23100
rect 16776 23032 16804 23072
rect 17865 23069 17877 23072
rect 17911 23100 17923 23103
rect 18782 23100 18788 23112
rect 17911 23072 18788 23100
rect 17911 23069 17923 23072
rect 17865 23063 17923 23069
rect 18782 23060 18788 23072
rect 18840 23060 18846 23112
rect 19150 23060 19156 23112
rect 19208 23100 19214 23112
rect 20165 23103 20223 23109
rect 20165 23100 20177 23103
rect 19208 23072 20177 23100
rect 19208 23060 19214 23072
rect 20165 23069 20177 23072
rect 20211 23069 20223 23103
rect 22922 23100 22928 23112
rect 20165 23063 20223 23069
rect 20272 23072 22928 23100
rect 15396 23004 16804 23032
rect 17681 23035 17739 23041
rect 17681 23001 17693 23035
rect 17727 23032 17739 23035
rect 17954 23032 17960 23044
rect 17727 23004 17960 23032
rect 17727 23001 17739 23004
rect 17681 22995 17739 23001
rect 17954 22992 17960 23004
rect 18012 22992 18018 23044
rect 18046 22992 18052 23044
rect 18104 23032 18110 23044
rect 20272 23032 20300 23072
rect 22922 23060 22928 23072
rect 22980 23060 22986 23112
rect 23290 23060 23296 23112
rect 23348 23100 23354 23112
rect 23860 23109 23888 23140
rect 24026 23128 24032 23140
rect 24084 23128 24090 23180
rect 24486 23168 24492 23180
rect 24447 23140 24492 23168
rect 24486 23128 24492 23140
rect 24544 23128 24550 23180
rect 23661 23103 23719 23109
rect 23661 23102 23673 23103
rect 23584 23100 23673 23102
rect 23348 23074 23673 23100
rect 23348 23072 23612 23074
rect 23348 23060 23354 23072
rect 23661 23069 23673 23074
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 23845 23103 23903 23109
rect 23845 23069 23857 23103
rect 23891 23069 23903 23103
rect 23845 23063 23903 23069
rect 24578 23060 24584 23112
rect 24636 23100 24642 23112
rect 24673 23103 24731 23109
rect 24673 23100 24685 23103
rect 24636 23072 24685 23100
rect 24636 23060 24642 23072
rect 24673 23069 24685 23072
rect 24719 23069 24731 23103
rect 24673 23063 24731 23069
rect 18104 23004 20300 23032
rect 20349 23035 20407 23041
rect 18104 22992 18110 23004
rect 20349 23001 20361 23035
rect 20395 23032 20407 23035
rect 20714 23032 20720 23044
rect 20395 23004 20720 23032
rect 20395 23001 20407 23004
rect 20349 22995 20407 23001
rect 13688 22936 14320 22964
rect 13688 22924 13694 22936
rect 14458 22924 14464 22976
rect 14516 22964 14522 22976
rect 20364 22964 20392 22995
rect 20714 22992 20720 23004
rect 20772 22992 20778 23044
rect 20806 22992 20812 23044
rect 20864 23032 20870 23044
rect 21085 23035 21143 23041
rect 21085 23032 21097 23035
rect 20864 23004 21097 23032
rect 20864 22992 20870 23004
rect 21085 23001 21097 23004
rect 21131 23032 21143 23035
rect 21726 23032 21732 23044
rect 21131 23004 21732 23032
rect 21131 23001 21143 23004
rect 21085 22995 21143 23001
rect 21726 22992 21732 23004
rect 21784 22992 21790 23044
rect 23753 23035 23811 23041
rect 23753 23001 23765 23035
rect 23799 23032 23811 23035
rect 24394 23032 24400 23044
rect 23799 23004 24400 23032
rect 23799 23001 23811 23004
rect 23753 22995 23811 23001
rect 24394 22992 24400 23004
rect 24452 22992 24458 23044
rect 24780 23032 24808 23208
rect 24857 23205 24869 23239
rect 24903 23205 24915 23239
rect 24857 23199 24915 23205
rect 24872 23100 24900 23199
rect 28074 23196 28080 23248
rect 28132 23236 28138 23248
rect 28132 23208 30328 23236
rect 28132 23196 28138 23208
rect 28902 23128 28908 23180
rect 28960 23168 28966 23180
rect 29086 23168 29092 23180
rect 28960 23140 29092 23168
rect 28960 23128 28966 23140
rect 29086 23128 29092 23140
rect 29144 23128 29150 23180
rect 25317 23103 25375 23109
rect 25317 23100 25329 23103
rect 24872 23072 25329 23100
rect 25317 23069 25329 23072
rect 25363 23069 25375 23103
rect 25317 23063 25375 23069
rect 28629 23103 28687 23109
rect 28629 23069 28641 23103
rect 28675 23100 28687 23103
rect 28994 23100 29000 23112
rect 28675 23072 29000 23100
rect 28675 23069 28687 23072
rect 28629 23063 28687 23069
rect 28994 23060 29000 23072
rect 29052 23060 29058 23112
rect 29822 23060 29828 23112
rect 29880 23100 29886 23112
rect 30116 23109 30236 23110
rect 30300 23109 30328 23208
rect 30116 23103 30251 23109
rect 30116 23100 30205 23103
rect 29880 23082 30205 23100
rect 29880 23072 30144 23082
rect 29880 23060 29886 23072
rect 30193 23069 30205 23082
rect 30239 23069 30251 23103
rect 30193 23063 30251 23069
rect 30282 23103 30340 23109
rect 30282 23069 30294 23103
rect 30328 23069 30340 23103
rect 30282 23063 30340 23069
rect 30374 23060 30380 23112
rect 30432 23100 30438 23112
rect 30561 23103 30619 23109
rect 30432 23072 30477 23100
rect 30432 23060 30438 23072
rect 30561 23069 30573 23103
rect 30607 23102 30619 23103
rect 30650 23102 30656 23112
rect 30607 23074 30656 23102
rect 30607 23069 30619 23074
rect 30561 23063 30619 23069
rect 30650 23060 30656 23074
rect 30708 23060 30714 23112
rect 31021 23103 31079 23109
rect 31021 23069 31033 23103
rect 31067 23100 31079 23103
rect 32490 23100 32496 23112
rect 31067 23072 32496 23100
rect 31067 23069 31079 23072
rect 31021 23063 31079 23069
rect 32490 23060 32496 23072
rect 32548 23060 32554 23112
rect 24780 23004 26924 23032
rect 21174 22964 21180 22976
rect 14516 22936 20392 22964
rect 21135 22936 21180 22964
rect 14516 22924 14522 22936
rect 21174 22924 21180 22936
rect 21232 22924 21238 22976
rect 23566 22924 23572 22976
rect 23624 22964 23630 22976
rect 24210 22964 24216 22976
rect 23624 22936 24216 22964
rect 23624 22924 23630 22936
rect 24210 22924 24216 22936
rect 24268 22924 24274 22976
rect 25501 22967 25559 22973
rect 25501 22933 25513 22967
rect 25547 22964 25559 22967
rect 26234 22964 26240 22976
rect 25547 22936 26240 22964
rect 25547 22933 25559 22936
rect 25501 22927 25559 22933
rect 26234 22924 26240 22936
rect 26292 22924 26298 22976
rect 26896 22964 26924 23004
rect 26970 22992 26976 23044
rect 27028 23032 27034 23044
rect 27246 23032 27252 23044
rect 27028 23004 27252 23032
rect 27028 22992 27034 23004
rect 27246 22992 27252 23004
rect 27304 23032 27310 23044
rect 28445 23035 28503 23041
rect 28445 23032 28457 23035
rect 27304 23004 28457 23032
rect 27304 22992 27310 23004
rect 28445 23001 28457 23004
rect 28491 23032 28503 23035
rect 29362 23032 29368 23044
rect 28491 23004 29368 23032
rect 28491 23001 28503 23004
rect 28445 22995 28503 23001
rect 29362 22992 29368 23004
rect 29420 22992 29426 23044
rect 30926 22964 30932 22976
rect 26896 22936 30932 22964
rect 30926 22924 30932 22936
rect 30984 22924 30990 22976
rect 31110 22964 31116 22976
rect 31071 22936 31116 22964
rect 31110 22924 31116 22936
rect 31168 22924 31174 22976
rect 1104 22874 48852 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 48852 22874
rect 1104 22800 48852 22822
rect 2590 22760 2596 22772
rect 2551 22732 2596 22760
rect 2590 22720 2596 22732
rect 2648 22720 2654 22772
rect 30558 22760 30564 22772
rect 2746 22732 28994 22760
rect 1486 22652 1492 22704
rect 1544 22692 1550 22704
rect 2746 22692 2774 22732
rect 12802 22692 12808 22704
rect 1544 22664 2774 22692
rect 12763 22664 12808 22692
rect 1544 22652 1550 22664
rect 12802 22652 12808 22664
rect 12860 22652 12866 22704
rect 13630 22692 13636 22704
rect 13591 22664 13636 22692
rect 13630 22652 13636 22664
rect 13688 22652 13694 22704
rect 14274 22692 14280 22704
rect 14187 22664 14280 22692
rect 14274 22652 14280 22664
rect 14332 22692 14338 22704
rect 14458 22692 14464 22704
rect 14332 22664 14464 22692
rect 14332 22652 14338 22664
rect 14458 22652 14464 22664
rect 14516 22652 14522 22704
rect 16945 22695 17003 22701
rect 16945 22661 16957 22695
rect 16991 22692 17003 22695
rect 17218 22692 17224 22704
rect 16991 22664 17224 22692
rect 16991 22661 17003 22664
rect 16945 22655 17003 22661
rect 17218 22652 17224 22664
rect 17276 22652 17282 22704
rect 17672 22695 17730 22701
rect 17672 22661 17684 22695
rect 17718 22692 17730 22695
rect 17862 22692 17868 22704
rect 17718 22664 17868 22692
rect 17718 22661 17730 22664
rect 17672 22655 17730 22661
rect 17862 22652 17868 22664
rect 17920 22652 17926 22704
rect 21174 22692 21180 22704
rect 19076 22664 21180 22692
rect 1854 22624 1860 22636
rect 1815 22596 1860 22624
rect 1854 22584 1860 22596
rect 1912 22584 1918 22636
rect 2498 22624 2504 22636
rect 2459 22596 2504 22624
rect 2498 22584 2504 22596
rect 2556 22584 2562 22636
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22593 12771 22627
rect 12713 22587 12771 22593
rect 12897 22627 12955 22633
rect 12897 22593 12909 22627
rect 12943 22624 12955 22627
rect 13262 22624 13268 22636
rect 12943 22596 13268 22624
rect 12943 22593 12955 22596
rect 12897 22587 12955 22593
rect 1946 22516 1952 22568
rect 2004 22556 2010 22568
rect 2590 22556 2596 22568
rect 2004 22528 2596 22556
rect 2004 22516 2010 22528
rect 2590 22516 2596 22528
rect 2648 22516 2654 22568
rect 12728 22488 12756 22587
rect 13262 22584 13268 22596
rect 13320 22584 13326 22636
rect 13354 22584 13360 22636
rect 13412 22624 13418 22636
rect 14090 22624 14096 22636
rect 13412 22596 13457 22624
rect 14051 22596 14096 22624
rect 13412 22584 13418 22596
rect 14090 22584 14096 22596
rect 14148 22584 14154 22636
rect 13170 22516 13176 22568
rect 13228 22556 13234 22568
rect 13446 22556 13452 22568
rect 13228 22528 13452 22556
rect 13228 22516 13234 22528
rect 13446 22516 13452 22528
rect 13504 22516 13510 22568
rect 13630 22556 13636 22568
rect 13591 22528 13636 22556
rect 13630 22516 13636 22528
rect 13688 22516 13694 22568
rect 14292 22556 14320 22652
rect 14366 22584 14372 22636
rect 14424 22624 14430 22636
rect 16761 22627 16819 22633
rect 14424 22596 14469 22624
rect 14424 22584 14430 22596
rect 16761 22593 16773 22627
rect 16807 22624 16819 22627
rect 19076 22624 19104 22664
rect 21174 22652 21180 22664
rect 21232 22652 21238 22704
rect 23842 22692 23848 22704
rect 23803 22664 23848 22692
rect 23842 22652 23848 22664
rect 23900 22652 23906 22704
rect 24670 22652 24676 22704
rect 24728 22692 24734 22704
rect 26145 22695 26203 22701
rect 24728 22664 25452 22692
rect 24728 22652 24734 22664
rect 16807 22596 19104 22624
rect 16807 22593 16819 22596
rect 16761 22587 16819 22593
rect 19150 22584 19156 22636
rect 19208 22624 19214 22636
rect 19521 22627 19579 22633
rect 19521 22624 19533 22627
rect 19208 22596 19533 22624
rect 19208 22584 19214 22596
rect 19521 22593 19533 22596
rect 19567 22624 19579 22627
rect 20533 22627 20591 22633
rect 20533 22624 20545 22627
rect 19567 22596 20545 22624
rect 19567 22593 19579 22596
rect 19521 22587 19579 22593
rect 20533 22593 20545 22596
rect 20579 22593 20591 22627
rect 20533 22587 20591 22593
rect 20717 22627 20775 22633
rect 20717 22593 20729 22627
rect 20763 22593 20775 22627
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 20717 22587 20775 22593
rect 13740 22528 14320 22556
rect 13740 22488 13768 22528
rect 15562 22516 15568 22568
rect 15620 22556 15626 22568
rect 17405 22559 17463 22565
rect 17405 22556 17417 22559
rect 15620 22528 17417 22556
rect 15620 22516 15626 22528
rect 17405 22525 17417 22528
rect 17451 22525 17463 22559
rect 19242 22556 19248 22568
rect 19203 22528 19248 22556
rect 17405 22519 17463 22525
rect 12728 22460 13768 22488
rect 14093 22491 14151 22497
rect 14093 22457 14105 22491
rect 14139 22488 14151 22491
rect 14550 22488 14556 22500
rect 14139 22460 14556 22488
rect 14139 22457 14151 22460
rect 14093 22451 14151 22457
rect 14550 22448 14556 22460
rect 14608 22448 14614 22500
rect 1946 22420 1952 22432
rect 1907 22392 1952 22420
rect 1946 22380 1952 22392
rect 2004 22380 2010 22432
rect 17420 22420 17448 22519
rect 19242 22516 19248 22528
rect 19300 22516 19306 22568
rect 18782 22488 18788 22500
rect 18743 22460 18788 22488
rect 18782 22448 18788 22460
rect 18840 22448 18846 22500
rect 20732 22488 20760 22587
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22094 22633 22100 22636
rect 22088 22587 22100 22633
rect 22152 22624 22158 22636
rect 22152 22596 22188 22624
rect 22094 22584 22100 22587
rect 22152 22584 22158 22596
rect 23014 22584 23020 22636
rect 23072 22624 23078 22636
rect 23753 22627 23811 22633
rect 23753 22624 23765 22627
rect 23072 22596 23765 22624
rect 23072 22584 23078 22596
rect 23753 22593 23765 22596
rect 23799 22624 23811 22627
rect 24578 22624 24584 22636
rect 23799 22596 24584 22624
rect 23799 22593 23811 22596
rect 23753 22587 23811 22593
rect 24578 22584 24584 22596
rect 24636 22584 24642 22636
rect 24854 22624 24860 22636
rect 24815 22596 24860 22624
rect 24854 22584 24860 22596
rect 24912 22584 24918 22636
rect 25130 22624 25136 22636
rect 25091 22596 25136 22624
rect 25130 22584 25136 22596
rect 25188 22584 25194 22636
rect 25424 22624 25452 22664
rect 26145 22661 26157 22695
rect 26191 22692 26203 22695
rect 26234 22692 26240 22704
rect 26191 22664 26240 22692
rect 26191 22661 26203 22664
rect 26145 22655 26203 22661
rect 26234 22652 26240 22664
rect 26292 22692 26298 22704
rect 26878 22692 26884 22704
rect 26292 22664 26884 22692
rect 26292 22652 26298 22664
rect 26878 22652 26884 22664
rect 26936 22652 26942 22704
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 25424 22596 26985 22624
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 27246 22624 27252 22636
rect 27207 22596 27252 22624
rect 26973 22587 27031 22593
rect 27246 22584 27252 22596
rect 27304 22584 27310 22636
rect 28966 22624 28994 22732
rect 29564 22732 30564 22760
rect 29319 22627 29377 22633
rect 29319 22624 29331 22627
rect 28966 22596 29331 22624
rect 29319 22593 29331 22596
rect 29365 22593 29377 22627
rect 29454 22624 29460 22636
rect 29415 22596 29460 22624
rect 29319 22587 29377 22593
rect 29454 22584 29460 22596
rect 29512 22584 29518 22636
rect 29564 22633 29592 22732
rect 30558 22720 30564 22732
rect 30616 22720 30622 22772
rect 30834 22720 30840 22772
rect 30892 22760 30898 22772
rect 31573 22763 31631 22769
rect 31573 22760 31585 22763
rect 30892 22732 31585 22760
rect 30892 22720 30898 22732
rect 31573 22729 31585 22732
rect 31619 22729 31631 22763
rect 31573 22723 31631 22729
rect 29822 22652 29828 22704
rect 29880 22692 29886 22704
rect 30852 22692 30880 22720
rect 46934 22692 46940 22704
rect 29880 22664 30880 22692
rect 34072 22664 46940 22692
rect 29880 22652 29886 22664
rect 29549 22627 29607 22633
rect 29549 22593 29561 22627
rect 29595 22593 29607 22627
rect 29730 22624 29736 22636
rect 29691 22596 29736 22624
rect 29549 22587 29607 22593
rect 29730 22584 29736 22596
rect 29788 22584 29794 22636
rect 30190 22624 30196 22636
rect 30151 22596 30196 22624
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 34072 22633 34100 22664
rect 46934 22652 46940 22664
rect 46992 22652 46998 22704
rect 30449 22627 30507 22633
rect 30449 22624 30461 22627
rect 30300 22596 30461 22624
rect 25041 22559 25099 22565
rect 25041 22525 25053 22559
rect 25087 22556 25099 22559
rect 25314 22556 25320 22568
rect 25087 22528 25320 22556
rect 25087 22525 25099 22528
rect 25041 22519 25099 22525
rect 25314 22516 25320 22528
rect 25372 22516 25378 22568
rect 30300 22556 30328 22596
rect 30449 22593 30461 22596
rect 30495 22593 30507 22627
rect 30449 22587 30507 22593
rect 34057 22627 34115 22633
rect 34057 22593 34069 22627
rect 34103 22593 34115 22627
rect 34057 22587 34115 22593
rect 34149 22627 34207 22633
rect 34149 22593 34161 22627
rect 34195 22593 34207 22627
rect 34149 22587 34207 22593
rect 34164 22556 34192 22587
rect 34238 22584 34244 22636
rect 34296 22624 34302 22636
rect 34425 22627 34483 22633
rect 34296 22596 34341 22624
rect 34296 22584 34302 22596
rect 34425 22593 34437 22627
rect 34471 22593 34483 22627
rect 48130 22624 48136 22636
rect 48091 22596 48136 22624
rect 34425 22587 34483 22593
rect 34440 22556 34468 22587
rect 48130 22584 48136 22596
rect 48188 22584 48194 22636
rect 30208 22528 30328 22556
rect 33704 22528 34192 22556
rect 34348 22528 34468 22556
rect 21358 22488 21364 22500
rect 20732 22460 21364 22488
rect 21358 22448 21364 22460
rect 21416 22488 21422 22500
rect 21416 22460 21864 22488
rect 21416 22448 21422 22460
rect 18690 22420 18696 22432
rect 17420 22392 18696 22420
rect 18690 22380 18696 22392
rect 18748 22380 18754 22432
rect 20901 22423 20959 22429
rect 20901 22389 20913 22423
rect 20947 22420 20959 22423
rect 21726 22420 21732 22432
rect 20947 22392 21732 22420
rect 20947 22389 20959 22392
rect 20901 22383 20959 22389
rect 21726 22380 21732 22392
rect 21784 22380 21790 22432
rect 21836 22420 21864 22460
rect 23934 22448 23940 22500
rect 23992 22488 23998 22500
rect 29089 22491 29147 22497
rect 23992 22460 25360 22488
rect 23992 22448 23998 22460
rect 23201 22423 23259 22429
rect 23201 22420 23213 22423
rect 21836 22392 23213 22420
rect 23201 22389 23213 22392
rect 23247 22389 23259 22423
rect 23201 22383 23259 22389
rect 25133 22423 25191 22429
rect 25133 22389 25145 22423
rect 25179 22420 25191 22423
rect 25222 22420 25228 22432
rect 25179 22392 25228 22420
rect 25179 22389 25191 22392
rect 25133 22383 25191 22389
rect 25222 22380 25228 22392
rect 25280 22380 25286 22432
rect 25332 22429 25360 22460
rect 29089 22457 29101 22491
rect 29135 22488 29147 22491
rect 30208 22488 30236 22528
rect 29135 22460 30236 22488
rect 29135 22457 29147 22460
rect 29089 22451 29147 22457
rect 25317 22423 25375 22429
rect 25317 22389 25329 22423
rect 25363 22389 25375 22423
rect 25317 22383 25375 22389
rect 25774 22380 25780 22432
rect 25832 22420 25838 22432
rect 26237 22423 26295 22429
rect 26237 22420 26249 22423
rect 25832 22392 26249 22420
rect 25832 22380 25838 22392
rect 26237 22389 26249 22392
rect 26283 22389 26295 22423
rect 26237 22383 26295 22389
rect 29454 22380 29460 22432
rect 29512 22420 29518 22432
rect 33704 22420 33732 22528
rect 29512 22392 33732 22420
rect 33781 22423 33839 22429
rect 29512 22380 29518 22392
rect 33781 22389 33793 22423
rect 33827 22420 33839 22423
rect 33870 22420 33876 22432
rect 33827 22392 33876 22420
rect 33827 22389 33839 22392
rect 33781 22383 33839 22389
rect 33870 22380 33876 22392
rect 33928 22380 33934 22432
rect 34072 22420 34100 22528
rect 34146 22448 34152 22500
rect 34204 22488 34210 22500
rect 34348 22488 34376 22528
rect 34204 22460 34376 22488
rect 34204 22448 34210 22460
rect 34514 22420 34520 22432
rect 34072 22392 34520 22420
rect 34514 22380 34520 22392
rect 34572 22380 34578 22432
rect 47578 22380 47584 22432
rect 47636 22420 47642 22432
rect 47949 22423 48007 22429
rect 47949 22420 47961 22423
rect 47636 22392 47961 22420
rect 47636 22380 47642 22392
rect 47949 22389 47961 22392
rect 47995 22389 48007 22423
rect 47949 22383 48007 22389
rect 1104 22330 48852 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 48852 22330
rect 1104 22256 48852 22278
rect 1946 22176 1952 22228
rect 2004 22216 2010 22228
rect 2004 22188 2774 22216
rect 2004 22176 2010 22188
rect 2746 22148 2774 22188
rect 13354 22176 13360 22228
rect 13412 22216 13418 22228
rect 14274 22216 14280 22228
rect 13412 22188 14280 22216
rect 13412 22176 13418 22188
rect 14274 22176 14280 22188
rect 14332 22176 14338 22228
rect 14384 22188 20668 22216
rect 14384 22148 14412 22188
rect 2746 22120 14412 22148
rect 14458 22108 14464 22160
rect 14516 22148 14522 22160
rect 20640 22148 20668 22188
rect 20714 22176 20720 22228
rect 20772 22216 20778 22228
rect 21818 22216 21824 22228
rect 20772 22188 21824 22216
rect 20772 22176 20778 22188
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 23661 22219 23719 22225
rect 23661 22185 23673 22219
rect 23707 22216 23719 22219
rect 23750 22216 23756 22228
rect 23707 22188 23756 22216
rect 23707 22185 23719 22188
rect 23661 22179 23719 22185
rect 23750 22176 23756 22188
rect 23808 22176 23814 22228
rect 24394 22216 24400 22228
rect 24355 22188 24400 22216
rect 24394 22176 24400 22188
rect 24452 22176 24458 22228
rect 24857 22219 24915 22225
rect 24857 22185 24869 22219
rect 24903 22216 24915 22219
rect 25130 22216 25136 22228
rect 24903 22188 25136 22216
rect 24903 22185 24915 22188
rect 24857 22179 24915 22185
rect 25130 22176 25136 22188
rect 25188 22176 25194 22228
rect 25498 22216 25504 22228
rect 25240 22188 25504 22216
rect 22278 22148 22284 22160
rect 14516 22120 14561 22148
rect 20640 22120 22284 22148
rect 14516 22108 14522 22120
rect 22278 22108 22284 22120
rect 22336 22108 22342 22160
rect 24486 22148 24492 22160
rect 23584 22120 24492 22148
rect 1670 22040 1676 22092
rect 1728 22080 1734 22092
rect 10873 22083 10931 22089
rect 10873 22080 10885 22083
rect 1728 22052 10885 22080
rect 1728 22040 1734 22052
rect 10873 22049 10885 22052
rect 10919 22080 10931 22083
rect 18046 22080 18052 22092
rect 10919 22052 18052 22080
rect 10919 22049 10931 22052
rect 10873 22043 10931 22049
rect 18046 22040 18052 22052
rect 18104 22040 18110 22092
rect 21910 22080 21916 22092
rect 21560 22052 21916 22080
rect 7006 21972 7012 22024
rect 7064 22012 7070 22024
rect 8202 22012 8208 22024
rect 7064 21984 8208 22012
rect 7064 21972 7070 21984
rect 8202 21972 8208 21984
rect 8260 22012 8266 22024
rect 9125 22015 9183 22021
rect 9125 22012 9137 22015
rect 8260 21984 9137 22012
rect 8260 21972 8266 21984
rect 9125 21981 9137 21984
rect 9171 21981 9183 22015
rect 10226 22012 10232 22024
rect 10187 21984 10232 22012
rect 9125 21975 9183 21981
rect 10226 21972 10232 21984
rect 10284 21972 10290 22024
rect 12986 21972 12992 22024
rect 13044 22012 13050 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13044 21984 14105 22012
rect 13044 21972 13050 21984
rect 14093 21981 14105 21984
rect 14139 22012 14151 22015
rect 14182 22012 14188 22024
rect 14139 21984 14188 22012
rect 14139 21981 14151 21984
rect 14093 21975 14151 21981
rect 14182 21972 14188 21984
rect 14240 21972 14246 22024
rect 14277 22015 14335 22021
rect 14277 21981 14289 22015
rect 14323 22012 14335 22015
rect 14366 22012 14372 22024
rect 14323 21984 14372 22012
rect 14323 21981 14335 21984
rect 14277 21975 14335 21981
rect 14366 21972 14372 21984
rect 14424 21972 14430 22024
rect 18279 22015 18337 22021
rect 18279 22012 18291 22015
rect 14476 21984 18291 22012
rect 8941 21947 8999 21953
rect 8941 21913 8953 21947
rect 8987 21944 8999 21947
rect 9214 21944 9220 21956
rect 8987 21916 9220 21944
rect 8987 21913 8999 21916
rect 8941 21907 8999 21913
rect 9214 21904 9220 21916
rect 9272 21904 9278 21956
rect 11057 21947 11115 21953
rect 11057 21913 11069 21947
rect 11103 21944 11115 21947
rect 11606 21944 11612 21956
rect 11103 21916 11612 21944
rect 11103 21913 11115 21916
rect 11057 21907 11115 21913
rect 11606 21904 11612 21916
rect 11664 21904 11670 21956
rect 12713 21947 12771 21953
rect 12713 21944 12725 21947
rect 12406 21916 12725 21944
rect 9309 21879 9367 21885
rect 9309 21845 9321 21879
rect 9355 21876 9367 21879
rect 9766 21876 9772 21888
rect 9355 21848 9772 21876
rect 9355 21845 9367 21848
rect 9309 21839 9367 21845
rect 9766 21836 9772 21848
rect 9824 21836 9830 21888
rect 10321 21879 10379 21885
rect 10321 21845 10333 21879
rect 10367 21876 10379 21879
rect 10594 21876 10600 21888
rect 10367 21848 10600 21876
rect 10367 21845 10379 21848
rect 10321 21839 10379 21845
rect 10594 21836 10600 21848
rect 10652 21836 10658 21888
rect 11238 21836 11244 21888
rect 11296 21876 11302 21888
rect 12406 21876 12434 21916
rect 12713 21913 12725 21916
rect 12759 21913 12771 21947
rect 12713 21907 12771 21913
rect 13078 21904 13084 21956
rect 13136 21944 13142 21956
rect 14476 21944 14504 21984
rect 18279 21981 18291 21984
rect 18325 21981 18337 22015
rect 18414 22012 18420 22024
rect 18375 21984 18420 22012
rect 18279 21975 18337 21981
rect 18414 21972 18420 21984
rect 18472 21972 18478 22024
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 18693 22015 18751 22021
rect 18564 21984 18609 22012
rect 18564 21972 18570 21984
rect 18693 21981 18705 22015
rect 18739 22012 18751 22015
rect 18782 22012 18788 22024
rect 18739 21984 18788 22012
rect 18739 21981 18751 21984
rect 18693 21975 18751 21981
rect 18782 21972 18788 21984
rect 18840 21972 18846 22024
rect 18874 21972 18880 22024
rect 18932 22012 18938 22024
rect 19245 22015 19303 22021
rect 19245 22012 19257 22015
rect 18932 21984 19257 22012
rect 18932 21972 18938 21984
rect 19245 21981 19257 21984
rect 19291 22012 19303 22015
rect 20714 22012 20720 22024
rect 19291 21984 20720 22012
rect 19291 21981 19303 21984
rect 19245 21975 19303 21981
rect 20714 21972 20720 21984
rect 20772 21972 20778 22024
rect 20990 21972 20996 22024
rect 21048 22012 21054 22024
rect 21560 22021 21588 22052
rect 21910 22040 21916 22052
rect 21968 22040 21974 22092
rect 21407 22015 21465 22021
rect 21407 22012 21419 22015
rect 21048 21984 21419 22012
rect 21048 21972 21054 21984
rect 21407 21981 21419 21984
rect 21453 21981 21465 22015
rect 21407 21975 21465 21981
rect 21542 22015 21600 22021
rect 21542 21981 21554 22015
rect 21588 21981 21600 22015
rect 21542 21975 21600 21981
rect 21637 22015 21695 22021
rect 21637 21981 21649 22015
rect 21683 22006 21695 22015
rect 21726 22006 21732 22024
rect 21683 21981 21732 22006
rect 21637 21978 21732 21981
rect 21637 21975 21695 21978
rect 21726 21972 21732 21978
rect 21784 21972 21790 22024
rect 21821 22015 21879 22021
rect 21821 21981 21833 22015
rect 21867 22012 21879 22015
rect 22646 22012 22652 22024
rect 21867 21984 22652 22012
rect 21867 21981 21879 21984
rect 21821 21975 21879 21981
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 23584 22012 23612 22120
rect 24486 22108 24492 22120
rect 24544 22108 24550 22160
rect 23952 22052 24716 22080
rect 23661 22015 23719 22021
rect 23661 22012 23673 22015
rect 23584 21984 23673 22012
rect 23661 21981 23673 21984
rect 23707 21981 23719 22015
rect 23842 22012 23848 22024
rect 23803 21984 23848 22012
rect 23661 21975 23719 21981
rect 23842 21972 23848 21984
rect 23900 21972 23906 22024
rect 13136 21916 14504 21944
rect 18049 21947 18107 21953
rect 13136 21904 13142 21916
rect 18049 21913 18061 21947
rect 18095 21944 18107 21947
rect 19490 21947 19548 21953
rect 19490 21944 19502 21947
rect 18095 21916 19502 21944
rect 18095 21913 18107 21916
rect 18049 21907 18107 21913
rect 19490 21913 19502 21916
rect 19536 21913 19548 21947
rect 19490 21907 19548 21913
rect 20254 21904 20260 21956
rect 20312 21944 20318 21956
rect 21177 21947 21235 21953
rect 21177 21944 21189 21947
rect 20312 21916 21189 21944
rect 20312 21904 20318 21916
rect 21177 21913 21189 21916
rect 21223 21913 21235 21947
rect 21177 21907 21235 21913
rect 23750 21904 23756 21956
rect 23808 21944 23814 21956
rect 23952 21944 23980 22052
rect 24688 22021 24716 22052
rect 25240 22024 25268 22188
rect 25498 22176 25504 22188
rect 25556 22176 25562 22228
rect 29730 22176 29736 22228
rect 29788 22216 29794 22228
rect 34146 22216 34152 22228
rect 29788 22188 34152 22216
rect 29788 22176 29794 22188
rect 34146 22176 34152 22188
rect 34204 22216 34210 22228
rect 34606 22216 34612 22228
rect 34204 22188 34612 22216
rect 34204 22176 34210 22188
rect 34606 22176 34612 22188
rect 34664 22176 34670 22228
rect 36630 22216 36636 22228
rect 34716 22188 36636 22216
rect 29086 22108 29092 22160
rect 29144 22148 29150 22160
rect 30650 22148 30656 22160
rect 29144 22120 30656 22148
rect 29144 22108 29150 22120
rect 30650 22108 30656 22120
rect 30708 22148 30714 22160
rect 32030 22148 32036 22160
rect 30708 22120 32036 22148
rect 30708 22108 30714 22120
rect 32030 22108 32036 22120
rect 32088 22108 32094 22160
rect 34238 22148 34244 22160
rect 33612 22120 34244 22148
rect 29733 22083 29791 22089
rect 29733 22049 29745 22083
rect 29779 22080 29791 22083
rect 31110 22080 31116 22092
rect 29779 22052 31116 22080
rect 29779 22049 29791 22052
rect 29733 22043 29791 22049
rect 31110 22040 31116 22052
rect 31168 22040 31174 22092
rect 33045 22083 33103 22089
rect 33045 22049 33057 22083
rect 33091 22080 33103 22083
rect 33612 22080 33640 22120
rect 34238 22108 34244 22120
rect 34296 22108 34302 22160
rect 34716 22080 34744 22188
rect 36630 22176 36636 22188
rect 36688 22176 36694 22228
rect 47762 22176 47768 22228
rect 47820 22216 47826 22228
rect 47857 22219 47915 22225
rect 47857 22216 47869 22219
rect 47820 22188 47869 22216
rect 47820 22176 47826 22188
rect 47857 22185 47869 22188
rect 47903 22185 47915 22219
rect 47857 22179 47915 22185
rect 47394 22080 47400 22092
rect 33091 22052 33640 22080
rect 33776 22052 34744 22080
rect 47355 22052 47400 22080
rect 33091 22049 33103 22052
rect 33045 22043 33103 22049
rect 24581 22015 24639 22021
rect 24581 21981 24593 22015
rect 24627 21981 24639 22015
rect 24581 21975 24639 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24394 21944 24400 21956
rect 23808 21916 23980 21944
rect 24355 21916 24400 21944
rect 23808 21904 23814 21916
rect 24394 21904 24400 21916
rect 24452 21904 24458 21956
rect 24596 21944 24624 21975
rect 25222 21972 25228 22024
rect 25280 21972 25286 22024
rect 25590 22012 25596 22024
rect 25551 21984 25596 22012
rect 25590 21972 25596 21984
rect 25648 22012 25654 22024
rect 27614 22012 27620 22024
rect 25648 21984 27620 22012
rect 25648 21972 25654 21984
rect 27614 21972 27620 21984
rect 27672 21972 27678 22024
rect 29546 22012 29552 22024
rect 29507 21984 29552 22012
rect 29546 21972 29552 21984
rect 29604 21972 29610 22024
rect 33776 22021 33804 22052
rect 47394 22040 47400 22052
rect 47452 22040 47458 22092
rect 33776 22015 33839 22021
rect 33776 21981 33793 22015
rect 33827 21981 33839 22015
rect 33781 21975 33839 21981
rect 33873 22015 33931 22021
rect 33873 21981 33885 22015
rect 33919 21981 33931 22015
rect 33873 21975 33931 21981
rect 24596 21916 24716 21944
rect 11296 21848 12434 21876
rect 11296 21836 11302 21848
rect 13446 21836 13452 21888
rect 13504 21876 13510 21888
rect 13630 21876 13636 21888
rect 13504 21848 13636 21876
rect 13504 21836 13510 21848
rect 13630 21836 13636 21848
rect 13688 21876 13694 21888
rect 14366 21876 14372 21888
rect 13688 21848 14372 21876
rect 13688 21836 13694 21848
rect 14366 21836 14372 21848
rect 14424 21876 14430 21888
rect 15838 21876 15844 21888
rect 14424 21848 15844 21876
rect 14424 21836 14430 21848
rect 15838 21836 15844 21848
rect 15896 21836 15902 21888
rect 20622 21876 20628 21888
rect 20583 21848 20628 21876
rect 20622 21836 20628 21848
rect 20680 21876 20686 21888
rect 24578 21876 24584 21888
rect 20680 21848 24584 21876
rect 20680 21836 20686 21848
rect 24578 21836 24584 21848
rect 24636 21836 24642 21888
rect 24688 21876 24716 21916
rect 25406 21904 25412 21956
rect 25464 21944 25470 21956
rect 25838 21947 25896 21953
rect 25838 21944 25850 21947
rect 25464 21916 25850 21944
rect 25464 21904 25470 21916
rect 25838 21913 25850 21916
rect 25884 21913 25896 21947
rect 27884 21947 27942 21953
rect 25838 21907 25896 21913
rect 25976 21916 27292 21944
rect 25976 21876 26004 21916
rect 24688 21848 26004 21876
rect 26973 21879 27031 21885
rect 26973 21845 26985 21879
rect 27019 21876 27031 21879
rect 27154 21876 27160 21888
rect 27019 21848 27160 21876
rect 27019 21845 27031 21848
rect 26973 21839 27031 21845
rect 27154 21836 27160 21848
rect 27212 21836 27218 21888
rect 27264 21876 27292 21916
rect 27884 21913 27896 21947
rect 27930 21944 27942 21947
rect 28258 21944 28264 21956
rect 27930 21916 28264 21944
rect 27930 21913 27942 21916
rect 27884 21907 27942 21913
rect 28258 21904 28264 21916
rect 28316 21904 28322 21956
rect 29914 21944 29920 21956
rect 28368 21916 29920 21944
rect 28368 21876 28396 21916
rect 29914 21904 29920 21916
rect 29972 21904 29978 21956
rect 31294 21904 31300 21956
rect 31352 21944 31358 21956
rect 31389 21947 31447 21953
rect 31389 21944 31401 21947
rect 31352 21916 31401 21944
rect 31352 21904 31358 21916
rect 31389 21913 31401 21916
rect 31435 21913 31447 21947
rect 32674 21944 32680 21956
rect 32635 21916 32680 21944
rect 31389 21907 31447 21913
rect 32674 21904 32680 21916
rect 32732 21904 32738 21956
rect 32858 21944 32864 21956
rect 32819 21916 32864 21944
rect 32858 21904 32864 21916
rect 32916 21904 32922 21956
rect 33888 21944 33916 21975
rect 33962 21972 33968 22024
rect 34020 22012 34026 22024
rect 34020 21984 34065 22012
rect 34020 21972 34026 21984
rect 34146 21972 34152 22024
rect 34204 22012 34210 22024
rect 34698 22012 34704 22024
rect 34204 21984 34249 22012
rect 34659 21984 34704 22012
rect 34204 21972 34210 21984
rect 34698 21972 34704 21984
rect 34756 21972 34762 22024
rect 47489 22015 47547 22021
rect 47489 21981 47501 22015
rect 47535 22012 47547 22015
rect 47578 22012 47584 22024
rect 47535 21984 47584 22012
rect 47535 21981 47547 21984
rect 47489 21975 47547 21981
rect 47578 21972 47584 21984
rect 47636 21972 47642 22024
rect 47854 22012 47860 22024
rect 47815 21984 47860 22012
rect 47854 21972 47860 21984
rect 47912 21972 47918 22024
rect 34514 21944 34520 21956
rect 33888 21916 34520 21944
rect 34514 21904 34520 21916
rect 34572 21904 34578 21956
rect 34946 21947 35004 21953
rect 34946 21913 34958 21947
rect 34992 21913 35004 21947
rect 34946 21907 35004 21913
rect 27264 21848 28396 21876
rect 28997 21879 29055 21885
rect 28997 21845 29009 21879
rect 29043 21876 29055 21879
rect 29546 21876 29552 21888
rect 29043 21848 29552 21876
rect 29043 21845 29055 21848
rect 28997 21839 29055 21845
rect 29546 21836 29552 21848
rect 29604 21836 29610 21888
rect 33505 21879 33563 21885
rect 33505 21845 33517 21879
rect 33551 21876 33563 21879
rect 34961 21876 34989 21907
rect 36078 21876 36084 21888
rect 33551 21848 34989 21876
rect 36039 21848 36084 21876
rect 33551 21845 33563 21848
rect 33505 21839 33563 21845
rect 36078 21836 36084 21848
rect 36136 21836 36142 21888
rect 36538 21836 36544 21888
rect 36596 21876 36602 21888
rect 48041 21879 48099 21885
rect 48041 21876 48053 21879
rect 36596 21848 48053 21876
rect 36596 21836 36602 21848
rect 48041 21845 48053 21848
rect 48087 21845 48099 21879
rect 48041 21839 48099 21845
rect 1104 21786 48852 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 48852 21786
rect 1104 21712 48852 21734
rect 8202 21632 8208 21684
rect 8260 21672 8266 21684
rect 8849 21675 8907 21681
rect 8849 21672 8861 21675
rect 8260 21644 8861 21672
rect 8260 21632 8266 21644
rect 8849 21641 8861 21644
rect 8895 21641 8907 21675
rect 11606 21672 11612 21684
rect 11567 21644 11612 21672
rect 8849 21635 8907 21641
rect 11606 21632 11612 21644
rect 11664 21632 11670 21684
rect 13449 21675 13507 21681
rect 13449 21641 13461 21675
rect 13495 21672 13507 21675
rect 13722 21672 13728 21684
rect 13495 21644 13728 21672
rect 13495 21641 13507 21644
rect 13449 21635 13507 21641
rect 13722 21632 13728 21644
rect 13780 21632 13786 21684
rect 18506 21632 18512 21684
rect 18564 21672 18570 21684
rect 19337 21675 19395 21681
rect 19337 21672 19349 21675
rect 18564 21644 19349 21672
rect 18564 21632 18570 21644
rect 19337 21641 19349 21644
rect 19383 21641 19395 21675
rect 26234 21672 26240 21684
rect 19337 21635 19395 21641
rect 20916 21644 26240 21672
rect 7736 21607 7794 21613
rect 7736 21573 7748 21607
rect 7782 21604 7794 21607
rect 9309 21607 9367 21613
rect 9309 21604 9321 21607
rect 7782 21576 9321 21604
rect 7782 21573 7794 21576
rect 7736 21567 7794 21573
rect 9309 21573 9321 21576
rect 9355 21573 9367 21607
rect 9309 21567 9367 21573
rect 9398 21564 9404 21616
rect 9456 21604 9462 21616
rect 19153 21607 19211 21613
rect 9456 21576 9720 21604
rect 9456 21564 9462 21576
rect 2406 21496 2412 21548
rect 2464 21536 2470 21548
rect 2464 21508 2774 21536
rect 2464 21496 2470 21508
rect 2746 21332 2774 21508
rect 9490 21496 9496 21548
rect 9548 21536 9554 21548
rect 9692 21545 9720 21576
rect 12406 21576 17080 21604
rect 9585 21539 9643 21545
rect 9585 21536 9597 21539
rect 9548 21508 9597 21536
rect 9548 21496 9554 21508
rect 9585 21505 9597 21508
rect 9631 21505 9643 21539
rect 9585 21499 9643 21505
rect 9677 21539 9735 21545
rect 9677 21505 9689 21539
rect 9723 21505 9735 21539
rect 9677 21499 9735 21505
rect 9766 21496 9772 21548
rect 9824 21536 9830 21548
rect 9953 21539 10011 21545
rect 9824 21508 9869 21536
rect 9824 21496 9830 21508
rect 9953 21505 9965 21539
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 7466 21468 7472 21480
rect 7427 21440 7472 21468
rect 7466 21428 7472 21440
rect 7524 21428 7530 21480
rect 9968 21468 9996 21499
rect 10226 21496 10232 21548
rect 10284 21536 10290 21548
rect 11517 21539 11575 21545
rect 11517 21536 11529 21539
rect 10284 21508 11529 21536
rect 10284 21496 10290 21508
rect 11517 21505 11529 21508
rect 11563 21536 11575 21539
rect 12406 21536 12434 21576
rect 12986 21536 12992 21548
rect 11563 21508 12434 21536
rect 12947 21508 12992 21536
rect 11563 21505 11575 21508
rect 11517 21499 11575 21505
rect 12986 21496 12992 21508
rect 13044 21496 13050 21548
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21536 13323 21539
rect 13354 21536 13360 21548
rect 13311 21508 13360 21536
rect 13311 21505 13323 21508
rect 13265 21499 13323 21505
rect 13354 21496 13360 21508
rect 13412 21496 13418 21548
rect 9646 21440 9996 21468
rect 13173 21471 13231 21477
rect 9490 21360 9496 21412
rect 9548 21400 9554 21412
rect 9646 21400 9674 21440
rect 13173 21437 13185 21471
rect 13219 21468 13231 21471
rect 14001 21471 14059 21477
rect 14001 21468 14013 21471
rect 13219 21440 14013 21468
rect 13219 21437 13231 21440
rect 13173 21431 13231 21437
rect 14001 21437 14013 21440
rect 14047 21437 14059 21471
rect 14274 21468 14280 21480
rect 14235 21440 14280 21468
rect 14001 21431 14059 21437
rect 9548 21372 9674 21400
rect 14016 21400 14044 21431
rect 14274 21428 14280 21440
rect 14332 21428 14338 21480
rect 17052 21468 17080 21576
rect 19153 21573 19165 21607
rect 19199 21604 19211 21607
rect 20622 21604 20628 21616
rect 19199 21576 20628 21604
rect 19199 21573 19211 21576
rect 19153 21567 19211 21573
rect 20622 21564 20628 21576
rect 20680 21564 20686 21616
rect 20717 21607 20775 21613
rect 20717 21573 20729 21607
rect 20763 21604 20775 21607
rect 20806 21604 20812 21616
rect 20763 21576 20812 21604
rect 20763 21573 20775 21576
rect 20717 21567 20775 21573
rect 20806 21564 20812 21576
rect 20864 21564 20870 21616
rect 17129 21539 17187 21545
rect 17129 21505 17141 21539
rect 17175 21536 17187 21539
rect 17862 21536 17868 21548
rect 17175 21508 17868 21536
rect 17175 21505 17187 21508
rect 17129 21499 17187 21505
rect 17862 21496 17868 21508
rect 17920 21496 17926 21548
rect 18969 21539 19027 21545
rect 18969 21505 18981 21539
rect 19015 21536 19027 21539
rect 19242 21536 19248 21548
rect 19015 21508 19248 21536
rect 19015 21505 19027 21508
rect 18969 21499 19027 21505
rect 19242 21496 19248 21508
rect 19300 21536 19306 21548
rect 19426 21536 19432 21548
rect 19300 21508 19432 21536
rect 19300 21496 19306 21508
rect 19426 21496 19432 21508
rect 19484 21496 19490 21548
rect 19981 21539 20039 21545
rect 19981 21505 19993 21539
rect 20027 21536 20039 21539
rect 20070 21536 20076 21548
rect 20027 21508 20076 21536
rect 20027 21505 20039 21508
rect 19981 21499 20039 21505
rect 20070 21496 20076 21508
rect 20128 21496 20134 21548
rect 20916 21468 20944 21644
rect 26234 21632 26240 21644
rect 26292 21632 26298 21684
rect 28258 21672 28264 21684
rect 26804 21644 27292 21672
rect 28219 21644 28264 21672
rect 20990 21564 20996 21616
rect 21048 21604 21054 21616
rect 21048 21576 26096 21604
rect 21048 21564 21054 21576
rect 21542 21496 21548 21548
rect 21600 21536 21606 21548
rect 22353 21539 22411 21545
rect 22353 21536 22365 21539
rect 21600 21508 22365 21536
rect 21600 21496 21606 21508
rect 22353 21505 22365 21508
rect 22399 21505 22411 21539
rect 22353 21499 22411 21505
rect 23658 21496 23664 21548
rect 23716 21536 23722 21548
rect 23937 21539 23995 21545
rect 23937 21536 23949 21539
rect 23716 21508 23949 21536
rect 23716 21496 23722 21508
rect 23937 21505 23949 21508
rect 23983 21505 23995 21539
rect 23937 21499 23995 21505
rect 24118 21496 24124 21548
rect 24176 21536 24182 21548
rect 25639 21539 25697 21545
rect 25639 21536 25651 21539
rect 24176 21508 25651 21536
rect 24176 21496 24182 21508
rect 25639 21505 25651 21508
rect 25685 21505 25697 21539
rect 25774 21536 25780 21548
rect 25735 21508 25780 21536
rect 25639 21499 25697 21505
rect 25774 21496 25780 21508
rect 25832 21496 25838 21548
rect 26068 21545 26096 21576
rect 26142 21564 26148 21616
rect 26200 21604 26206 21616
rect 26804 21604 26832 21644
rect 26970 21604 26976 21616
rect 26200 21576 26832 21604
rect 26931 21576 26976 21604
rect 26200 21564 26206 21576
rect 26970 21564 26976 21576
rect 27028 21564 27034 21616
rect 25869 21539 25927 21545
rect 25869 21505 25881 21539
rect 25915 21505 25927 21539
rect 25869 21499 25927 21505
rect 26053 21539 26111 21545
rect 26053 21505 26065 21539
rect 26099 21505 26111 21539
rect 27154 21536 27160 21548
rect 27115 21508 27160 21536
rect 26053 21499 26111 21505
rect 17052 21440 20944 21468
rect 21174 21428 21180 21480
rect 21232 21468 21238 21480
rect 21818 21468 21824 21480
rect 21232 21440 21824 21468
rect 21232 21428 21238 21440
rect 21818 21428 21824 21440
rect 21876 21468 21882 21480
rect 22097 21471 22155 21477
rect 22097 21468 22109 21471
rect 21876 21440 22109 21468
rect 21876 21428 21882 21440
rect 22097 21437 22109 21440
rect 22143 21437 22155 21471
rect 22097 21431 22155 21437
rect 24026 21428 24032 21480
rect 24084 21468 24090 21480
rect 24762 21468 24768 21480
rect 24084 21440 24768 21468
rect 24084 21428 24090 21440
rect 24762 21428 24768 21440
rect 24820 21428 24826 21480
rect 25406 21468 25412 21480
rect 25367 21440 25412 21468
rect 25406 21428 25412 21440
rect 25464 21428 25470 21480
rect 25884 21468 25912 21499
rect 27154 21496 27160 21508
rect 27212 21496 27218 21548
rect 27264 21536 27292 21644
rect 28258 21632 28264 21644
rect 28316 21632 28322 21684
rect 30558 21672 30564 21684
rect 30519 21644 30564 21672
rect 30558 21632 30564 21644
rect 30616 21632 30622 21684
rect 47762 21672 47768 21684
rect 30668 21644 47768 21672
rect 29178 21604 29184 21616
rect 28506 21576 29184 21604
rect 28506 21545 28534 21576
rect 29178 21564 29184 21576
rect 29236 21564 29242 21616
rect 29362 21604 29368 21616
rect 29323 21576 29368 21604
rect 29362 21564 29368 21576
rect 29420 21564 29426 21616
rect 29546 21604 29552 21616
rect 29507 21576 29552 21604
rect 29546 21564 29552 21576
rect 29604 21564 29610 21616
rect 29638 21564 29644 21616
rect 29696 21604 29702 21616
rect 30668 21604 30696 21644
rect 47762 21632 47768 21644
rect 47820 21632 47826 21684
rect 34698 21604 34704 21616
rect 29696 21576 30696 21604
rect 33796 21576 34704 21604
rect 29696 21564 29702 21576
rect 28491 21539 28549 21545
rect 28491 21536 28503 21539
rect 27264 21508 28503 21536
rect 28491 21505 28503 21508
rect 28537 21505 28549 21539
rect 28491 21499 28549 21505
rect 28629 21539 28687 21545
rect 28629 21505 28641 21539
rect 28675 21505 28687 21539
rect 28629 21499 28687 21505
rect 28721 21539 28779 21545
rect 28721 21505 28733 21539
rect 28767 21505 28779 21539
rect 28902 21536 28908 21548
rect 28863 21508 28908 21536
rect 28721 21499 28779 21505
rect 27341 21471 27399 21477
rect 27341 21468 27353 21471
rect 25884 21440 27353 21468
rect 27341 21437 27353 21440
rect 27387 21437 27399 21471
rect 27341 21431 27399 21437
rect 28074 21428 28080 21480
rect 28132 21468 28138 21480
rect 28644 21468 28672 21499
rect 28132 21440 28672 21468
rect 28736 21468 28764 21499
rect 28902 21496 28908 21508
rect 28960 21496 28966 21548
rect 30193 21539 30251 21545
rect 30193 21536 30205 21539
rect 30188 21505 30205 21536
rect 30239 21505 30251 21539
rect 30188 21499 30251 21505
rect 30377 21539 30435 21545
rect 30377 21505 30389 21539
rect 30423 21536 30435 21539
rect 30834 21536 30840 21548
rect 30423 21508 30840 21536
rect 30423 21505 30435 21508
rect 30377 21499 30435 21505
rect 29733 21471 29791 21477
rect 29733 21468 29745 21471
rect 28736 21440 29745 21468
rect 28132 21428 28138 21440
rect 29733 21437 29745 21440
rect 29779 21437 29791 21471
rect 29733 21431 29791 21437
rect 30188 21468 30216 21499
rect 30834 21496 30840 21508
rect 30892 21496 30898 21548
rect 33796 21545 33824 21576
rect 34698 21564 34704 21576
rect 34756 21564 34762 21616
rect 47946 21604 47952 21616
rect 47907 21576 47952 21604
rect 47946 21564 47952 21576
rect 48004 21564 48010 21616
rect 33781 21539 33839 21545
rect 33781 21505 33793 21539
rect 33827 21505 33839 21539
rect 33781 21499 33839 21505
rect 33870 21496 33876 21548
rect 33928 21536 33934 21548
rect 34037 21539 34095 21545
rect 34037 21536 34049 21539
rect 33928 21508 34049 21536
rect 33928 21496 33934 21508
rect 34037 21505 34049 21508
rect 34083 21505 34095 21539
rect 34037 21499 34095 21505
rect 32674 21468 32680 21480
rect 30188 21440 32680 21468
rect 15654 21400 15660 21412
rect 14016 21372 15660 21400
rect 9548 21360 9554 21372
rect 15654 21360 15660 21372
rect 15712 21360 15718 21412
rect 17310 21400 17316 21412
rect 17271 21372 17316 21400
rect 17310 21360 17316 21372
rect 17368 21360 17374 21412
rect 18414 21360 18420 21412
rect 18472 21400 18478 21412
rect 19242 21400 19248 21412
rect 18472 21372 19248 21400
rect 18472 21360 18478 21372
rect 19242 21360 19248 21372
rect 19300 21400 19306 21412
rect 20901 21403 20959 21409
rect 20901 21400 20913 21403
rect 19300 21372 20913 21400
rect 19300 21360 19306 21372
rect 20901 21369 20913 21372
rect 20947 21369 20959 21403
rect 20901 21363 20959 21369
rect 24578 21360 24584 21412
rect 24636 21400 24642 21412
rect 29638 21400 29644 21412
rect 24636 21372 29644 21400
rect 24636 21360 24642 21372
rect 29638 21360 29644 21372
rect 29696 21360 29702 21412
rect 13078 21332 13084 21344
rect 2746 21304 13084 21332
rect 13078 21292 13084 21304
rect 13136 21292 13142 21344
rect 13265 21335 13323 21341
rect 13265 21301 13277 21335
rect 13311 21332 13323 21335
rect 13446 21332 13452 21344
rect 13311 21304 13452 21332
rect 13311 21301 13323 21304
rect 13265 21295 13323 21301
rect 13446 21292 13452 21304
rect 13504 21292 13510 21344
rect 13998 21292 14004 21344
rect 14056 21332 14062 21344
rect 17494 21332 17500 21344
rect 14056 21304 17500 21332
rect 14056 21292 14062 21304
rect 17494 21292 17500 21304
rect 17552 21332 17558 21344
rect 17957 21335 18015 21341
rect 17957 21332 17969 21335
rect 17552 21304 17969 21332
rect 17552 21292 17558 21304
rect 17957 21301 17969 21304
rect 18003 21301 18015 21335
rect 17957 21295 18015 21301
rect 19426 21292 19432 21344
rect 19484 21332 19490 21344
rect 19797 21335 19855 21341
rect 19797 21332 19809 21335
rect 19484 21304 19809 21332
rect 19484 21292 19490 21304
rect 19797 21301 19809 21304
rect 19843 21301 19855 21335
rect 19797 21295 19855 21301
rect 23474 21292 23480 21344
rect 23532 21332 23538 21344
rect 24167 21335 24225 21341
rect 23532 21304 23577 21332
rect 23532 21292 23538 21304
rect 24167 21301 24179 21335
rect 24213 21332 24225 21335
rect 24486 21332 24492 21344
rect 24213 21304 24492 21332
rect 24213 21301 24225 21304
rect 24167 21295 24225 21301
rect 24486 21292 24492 21304
rect 24544 21332 24550 21344
rect 30188 21332 30216 21440
rect 32674 21428 32680 21440
rect 32732 21428 32738 21480
rect 24544 21304 30216 21332
rect 24544 21292 24550 21304
rect 31846 21292 31852 21344
rect 31904 21332 31910 21344
rect 32858 21332 32864 21344
rect 31904 21304 32864 21332
rect 31904 21292 31910 21304
rect 32858 21292 32864 21304
rect 32916 21332 32922 21344
rect 35161 21335 35219 21341
rect 35161 21332 35173 21335
rect 32916 21304 35173 21332
rect 32916 21292 32922 21304
rect 35161 21301 35173 21304
rect 35207 21301 35219 21335
rect 48038 21332 48044 21344
rect 47999 21304 48044 21332
rect 35161 21295 35219 21301
rect 48038 21292 48044 21304
rect 48096 21292 48102 21344
rect 1104 21242 48852 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 48852 21242
rect 1104 21168 48852 21190
rect 4614 21088 4620 21140
rect 4672 21128 4678 21140
rect 4672 21100 17172 21128
rect 4672 21088 4678 21100
rect 3970 21020 3976 21072
rect 4028 21060 4034 21072
rect 15654 21060 15660 21072
rect 4028 21032 11100 21060
rect 15615 21032 15660 21060
rect 4028 21020 4034 21032
rect 4062 20952 4068 21004
rect 4120 20992 4126 21004
rect 6917 20995 6975 21001
rect 6917 20992 6929 20995
rect 4120 20964 6929 20992
rect 4120 20952 4126 20964
rect 6917 20961 6929 20964
rect 6963 20961 6975 20995
rect 10594 20992 10600 21004
rect 10555 20964 10600 20992
rect 6917 20955 6975 20961
rect 10594 20952 10600 20964
rect 10652 20952 10658 21004
rect 11072 21001 11100 21032
rect 15654 21020 15660 21032
rect 15712 21020 15718 21072
rect 11057 20995 11115 21001
rect 11057 20961 11069 20995
rect 11103 20961 11115 20995
rect 11057 20955 11115 20961
rect 6273 20927 6331 20933
rect 6273 20893 6285 20927
rect 6319 20893 6331 20927
rect 6273 20887 6331 20893
rect 6288 20788 6316 20887
rect 9030 20884 9036 20936
rect 9088 20924 9094 20936
rect 9171 20927 9229 20933
rect 9171 20924 9183 20927
rect 9088 20896 9183 20924
rect 9088 20884 9094 20896
rect 9171 20893 9183 20896
rect 9217 20893 9229 20927
rect 9303 20921 9309 20933
rect 9264 20893 9309 20921
rect 9171 20887 9229 20893
rect 9303 20881 9309 20893
rect 9361 20881 9367 20933
rect 9398 20884 9404 20936
rect 9456 20924 9462 20936
rect 9585 20927 9643 20933
rect 9456 20896 9501 20924
rect 9456 20884 9462 20896
rect 9585 20893 9597 20927
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 10413 20927 10471 20933
rect 10413 20893 10425 20927
rect 10459 20893 10471 20927
rect 10413 20887 10471 20893
rect 6454 20856 6460 20868
rect 6415 20828 6460 20856
rect 6454 20816 6460 20828
rect 6512 20816 6518 20868
rect 9600 20856 9628 20887
rect 9508 20828 9628 20856
rect 10428 20856 10456 20887
rect 13170 20884 13176 20936
rect 13228 20924 13234 20936
rect 14277 20927 14335 20933
rect 14277 20924 14289 20927
rect 13228 20896 14289 20924
rect 13228 20884 13234 20896
rect 14277 20893 14289 20896
rect 14323 20893 14335 20927
rect 14277 20887 14335 20893
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20924 16175 20927
rect 16163 20896 16528 20924
rect 16163 20893 16175 20896
rect 16117 20887 16175 20893
rect 16500 20868 16528 20896
rect 10778 20856 10784 20868
rect 10428 20828 10784 20856
rect 9508 20800 9536 20828
rect 10778 20816 10784 20828
rect 10836 20816 10842 20868
rect 14550 20865 14556 20868
rect 14544 20819 14556 20865
rect 14608 20856 14614 20868
rect 16384 20859 16442 20865
rect 14608 20828 14644 20856
rect 14550 20816 14556 20819
rect 14608 20816 14614 20828
rect 16384 20825 16396 20859
rect 16430 20825 16442 20859
rect 16384 20819 16442 20825
rect 8202 20788 8208 20800
rect 6288 20760 8208 20788
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 8938 20788 8944 20800
rect 8899 20760 8944 20788
rect 8938 20748 8944 20760
rect 8996 20748 9002 20800
rect 9490 20748 9496 20800
rect 9548 20748 9554 20800
rect 16408 20788 16436 20819
rect 16482 20816 16488 20868
rect 16540 20816 16546 20868
rect 17144 20856 17172 21100
rect 18690 21088 18696 21140
rect 18748 21128 18754 21140
rect 20990 21128 20996 21140
rect 18748 21100 20996 21128
rect 18748 21088 18754 21100
rect 20990 21088 20996 21100
rect 21048 21088 21054 21140
rect 21100 21100 21833 21128
rect 20901 21063 20959 21069
rect 20901 21029 20913 21063
rect 20947 21060 20959 21063
rect 21100 21060 21128 21100
rect 20947 21032 21128 21060
rect 21361 21063 21419 21069
rect 20947 21029 20959 21032
rect 20901 21023 20959 21029
rect 21361 21029 21373 21063
rect 21407 21060 21419 21063
rect 21542 21060 21548 21072
rect 21407 21032 21548 21060
rect 21407 21029 21419 21032
rect 21361 21023 21419 21029
rect 21542 21020 21548 21032
rect 21600 21020 21606 21072
rect 17862 20952 17868 21004
rect 17920 20992 17926 21004
rect 21450 20992 21456 21004
rect 17920 20964 21456 20992
rect 17920 20952 17926 20964
rect 19720 20933 19748 20964
rect 21450 20952 21456 20964
rect 21508 20952 21514 21004
rect 21652 20992 21680 21100
rect 21805 21060 21833 21100
rect 25130 21088 25136 21140
rect 25188 21128 25194 21140
rect 33962 21128 33968 21140
rect 25188 21100 33824 21128
rect 33923 21100 33968 21128
rect 25188 21088 25194 21100
rect 29454 21060 29460 21072
rect 21805 21032 29460 21060
rect 29454 21020 29460 21032
rect 29512 21020 29518 21072
rect 31110 21020 31116 21072
rect 31168 21060 31174 21072
rect 33796 21060 33824 21100
rect 33962 21088 33968 21100
rect 34020 21088 34026 21140
rect 36538 21060 36544 21072
rect 31168 21032 33732 21060
rect 33796 21032 36544 21060
rect 31168 21020 31174 21032
rect 24765 20995 24823 21001
rect 24765 20992 24777 20995
rect 21652 20964 21772 20992
rect 19705 20927 19763 20933
rect 19705 20893 19717 20927
rect 19751 20893 19763 20927
rect 20714 20924 20720 20936
rect 20675 20896 20720 20924
rect 19705 20887 19763 20893
rect 20714 20884 20720 20896
rect 20772 20884 20778 20936
rect 21637 20927 21695 20933
rect 21744 20927 21772 20964
rect 21928 20964 24777 20992
rect 21842 20927 21900 20933
rect 21637 20924 21649 20927
rect 20815 20896 21649 20924
rect 20815 20856 20843 20896
rect 21637 20893 21649 20896
rect 21683 20893 21695 20927
rect 21637 20887 21695 20893
rect 21742 20921 21800 20927
rect 21742 20887 21754 20921
rect 21788 20887 21800 20921
rect 21842 20893 21854 20927
rect 21888 20924 21900 20927
rect 21928 20924 21956 20964
rect 24765 20961 24777 20964
rect 24811 20961 24823 20995
rect 24765 20955 24823 20961
rect 26881 20995 26939 21001
rect 26881 20961 26893 20995
rect 26927 20992 26939 20995
rect 27154 20992 27160 21004
rect 26927 20964 27160 20992
rect 26927 20961 26939 20964
rect 26881 20955 26939 20961
rect 27154 20952 27160 20964
rect 27212 20952 27218 21004
rect 33704 20992 33732 21032
rect 36538 21020 36544 21032
rect 36596 21020 36602 21072
rect 33704 20964 33824 20992
rect 21888 20896 21956 20924
rect 22005 20927 22063 20933
rect 21888 20893 21900 20896
rect 21842 20887 21900 20893
rect 22005 20893 22017 20927
rect 22051 20924 22063 20927
rect 22094 20924 22100 20936
rect 22051 20896 22100 20924
rect 22051 20893 22063 20896
rect 22005 20887 22063 20893
rect 21742 20881 21800 20887
rect 22094 20884 22100 20896
rect 22152 20884 22158 20936
rect 23474 20884 23480 20936
rect 23532 20924 23538 20936
rect 24397 20927 24455 20933
rect 23532 20896 24348 20924
rect 23532 20884 23538 20896
rect 22557 20859 22615 20865
rect 22557 20856 22569 20859
rect 17144 20828 20843 20856
rect 21928 20828 22569 20856
rect 16758 20788 16764 20800
rect 16408 20760 16764 20788
rect 16758 20748 16764 20760
rect 16816 20748 16822 20800
rect 16850 20748 16856 20800
rect 16908 20788 16914 20800
rect 17497 20791 17555 20797
rect 17497 20788 17509 20791
rect 16908 20760 17509 20788
rect 16908 20748 16914 20760
rect 17497 20757 17509 20760
rect 17543 20757 17555 20791
rect 17497 20751 17555 20757
rect 18782 20748 18788 20800
rect 18840 20788 18846 20800
rect 19797 20791 19855 20797
rect 19797 20788 19809 20791
rect 18840 20760 19809 20788
rect 18840 20748 18846 20760
rect 19797 20757 19809 20760
rect 19843 20788 19855 20791
rect 20990 20788 20996 20800
rect 19843 20760 20996 20788
rect 19843 20757 19855 20760
rect 19797 20751 19855 20757
rect 20990 20748 20996 20760
rect 21048 20748 21054 20800
rect 21450 20748 21456 20800
rect 21508 20788 21514 20800
rect 21928 20788 21956 20828
rect 22557 20825 22569 20828
rect 22603 20856 22615 20859
rect 23661 20859 23719 20865
rect 22603 20828 22784 20856
rect 22603 20825 22615 20828
rect 22557 20819 22615 20825
rect 22646 20788 22652 20800
rect 21508 20760 21956 20788
rect 22607 20760 22652 20788
rect 21508 20748 21514 20760
rect 22646 20748 22652 20760
rect 22704 20748 22710 20800
rect 22756 20788 22784 20828
rect 23661 20825 23673 20859
rect 23707 20856 23719 20859
rect 24026 20856 24032 20868
rect 23707 20828 24032 20856
rect 23707 20825 23719 20828
rect 23661 20819 23719 20825
rect 24026 20816 24032 20828
rect 24084 20816 24090 20868
rect 24320 20856 24348 20896
rect 24397 20893 24409 20927
rect 24443 20924 24455 20927
rect 24486 20924 24492 20936
rect 24443 20896 24492 20924
rect 24443 20893 24455 20896
rect 24397 20887 24455 20893
rect 24486 20884 24492 20896
rect 24544 20884 24550 20936
rect 26234 20924 26240 20936
rect 26195 20896 26240 20924
rect 26234 20884 26240 20896
rect 26292 20884 26298 20936
rect 31202 20884 31208 20936
rect 31260 20924 31266 20936
rect 31527 20927 31585 20933
rect 31527 20924 31539 20927
rect 31260 20896 31539 20924
rect 31260 20884 31266 20896
rect 31527 20893 31539 20896
rect 31573 20893 31585 20927
rect 31527 20887 31585 20893
rect 31665 20927 31723 20933
rect 31665 20893 31677 20927
rect 31711 20893 31723 20927
rect 31665 20887 31723 20893
rect 31778 20924 31836 20930
rect 31778 20890 31790 20924
rect 31824 20921 31836 20924
rect 31941 20927 31999 20933
rect 31824 20893 31892 20921
rect 31824 20890 31836 20893
rect 24581 20859 24639 20865
rect 24581 20856 24593 20859
rect 24320 20828 24593 20856
rect 24581 20825 24593 20828
rect 24627 20856 24639 20859
rect 26142 20856 26148 20868
rect 24627 20828 26148 20856
rect 24627 20825 24639 20828
rect 24581 20819 24639 20825
rect 26142 20816 26148 20828
rect 26200 20816 26206 20868
rect 26329 20859 26387 20865
rect 26329 20825 26341 20859
rect 26375 20856 26387 20859
rect 27065 20859 27123 20865
rect 27065 20856 27077 20859
rect 26375 20828 27077 20856
rect 26375 20825 26387 20828
rect 26329 20819 26387 20825
rect 27065 20825 27077 20828
rect 27111 20825 27123 20859
rect 28718 20856 28724 20868
rect 28679 20828 28724 20856
rect 27065 20819 27123 20825
rect 28718 20816 28724 20828
rect 28776 20816 28782 20868
rect 30650 20816 30656 20868
rect 30708 20856 30714 20868
rect 31680 20856 31708 20887
rect 31778 20884 31836 20890
rect 30708 20828 31708 20856
rect 31864 20856 31892 20893
rect 31941 20893 31953 20927
rect 31987 20924 31999 20927
rect 32030 20924 32036 20936
rect 31987 20896 32036 20924
rect 31987 20893 31999 20896
rect 31941 20887 31999 20893
rect 32030 20884 32036 20896
rect 32088 20884 32094 20936
rect 32582 20924 32588 20936
rect 32543 20896 32588 20924
rect 32582 20884 32588 20896
rect 32640 20884 32646 20936
rect 32674 20884 32680 20936
rect 32732 20924 32738 20936
rect 33597 20927 33655 20933
rect 33597 20924 33609 20927
rect 32732 20896 33609 20924
rect 32732 20884 32738 20896
rect 33597 20893 33609 20896
rect 33643 20924 33655 20927
rect 33686 20924 33692 20936
rect 33643 20896 33692 20924
rect 33643 20893 33655 20896
rect 33597 20887 33655 20893
rect 33686 20884 33692 20896
rect 33744 20884 33750 20936
rect 33796 20933 33824 20964
rect 33781 20927 33839 20933
rect 33781 20893 33793 20927
rect 33827 20924 33839 20927
rect 36078 20924 36084 20936
rect 33827 20896 36084 20924
rect 33827 20893 33839 20896
rect 33781 20887 33839 20893
rect 36078 20884 36084 20896
rect 36136 20884 36142 20936
rect 31864 20828 32260 20856
rect 30708 20816 30714 20828
rect 23753 20791 23811 20797
rect 23753 20788 23765 20791
rect 22756 20760 23765 20788
rect 23753 20757 23765 20760
rect 23799 20788 23811 20791
rect 27982 20788 27988 20800
rect 23799 20760 27988 20788
rect 23799 20757 23811 20760
rect 23753 20751 23811 20757
rect 27982 20748 27988 20760
rect 28040 20748 28046 20800
rect 31297 20791 31355 20797
rect 31297 20757 31309 20791
rect 31343 20788 31355 20791
rect 32122 20788 32128 20800
rect 31343 20760 32128 20788
rect 31343 20757 31355 20760
rect 31297 20751 31355 20757
rect 32122 20748 32128 20760
rect 32180 20748 32186 20800
rect 32232 20788 32260 20828
rect 32306 20816 32312 20868
rect 32364 20856 32370 20868
rect 32401 20859 32459 20865
rect 32401 20856 32413 20859
rect 32364 20828 32413 20856
rect 32364 20816 32370 20828
rect 32401 20825 32413 20828
rect 32447 20825 32459 20859
rect 32401 20819 32459 20825
rect 32769 20791 32827 20797
rect 32769 20788 32781 20791
rect 32232 20760 32781 20788
rect 32769 20757 32781 20760
rect 32815 20757 32827 20791
rect 32769 20751 32827 20757
rect 1104 20698 48852 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 48852 20698
rect 1104 20624 48852 20646
rect 6454 20584 6460 20596
rect 6415 20556 6460 20584
rect 6454 20544 6460 20556
rect 6512 20544 6518 20596
rect 8202 20544 8208 20596
rect 8260 20584 8266 20596
rect 8757 20587 8815 20593
rect 8757 20584 8769 20587
rect 8260 20556 8769 20584
rect 8260 20544 8266 20556
rect 8757 20553 8769 20556
rect 8803 20553 8815 20587
rect 8757 20547 8815 20553
rect 7466 20516 7472 20528
rect 7379 20488 7472 20516
rect 6362 20448 6368 20460
rect 6323 20420 6368 20448
rect 6362 20408 6368 20420
rect 6420 20408 6426 20460
rect 7392 20457 7420 20488
rect 7466 20476 7472 20488
rect 7524 20516 7530 20528
rect 7834 20516 7840 20528
rect 7524 20488 7840 20516
rect 7524 20476 7530 20488
rect 7834 20476 7840 20488
rect 7892 20476 7898 20528
rect 8772 20516 8800 20547
rect 9398 20544 9404 20596
rect 9456 20584 9462 20596
rect 9585 20587 9643 20593
rect 9585 20584 9597 20587
rect 9456 20556 9597 20584
rect 9456 20544 9462 20556
rect 9585 20553 9597 20556
rect 9631 20553 9643 20587
rect 9585 20547 9643 20553
rect 14461 20587 14519 20593
rect 14461 20553 14473 20587
rect 14507 20584 14519 20587
rect 14550 20584 14556 20596
rect 14507 20556 14556 20584
rect 14507 20553 14519 20556
rect 14461 20547 14519 20553
rect 14550 20544 14556 20556
rect 14608 20544 14614 20596
rect 16669 20587 16727 20593
rect 16669 20553 16681 20587
rect 16715 20584 16727 20587
rect 16758 20584 16764 20596
rect 16715 20556 16764 20584
rect 16715 20553 16727 20556
rect 16669 20547 16727 20553
rect 16758 20544 16764 20556
rect 16816 20544 16822 20596
rect 23474 20584 23480 20596
rect 16868 20556 23480 20584
rect 16868 20516 16896 20556
rect 23474 20544 23480 20556
rect 23532 20544 23538 20596
rect 23768 20556 41414 20584
rect 17678 20516 17684 20528
rect 8772 20488 9444 20516
rect 7377 20451 7435 20457
rect 7377 20417 7389 20451
rect 7423 20417 7435 20451
rect 7377 20411 7435 20417
rect 7644 20451 7702 20457
rect 7644 20417 7656 20451
rect 7690 20448 7702 20451
rect 8938 20448 8944 20460
rect 7690 20420 8944 20448
rect 7690 20417 7702 20420
rect 7644 20411 7702 20417
rect 8938 20408 8944 20420
rect 8996 20408 9002 20460
rect 9214 20448 9220 20460
rect 9175 20420 9220 20448
rect 9214 20408 9220 20420
rect 9272 20408 9278 20460
rect 9416 20457 9444 20488
rect 14752 20488 16896 20516
rect 16940 20488 17684 20516
rect 9401 20451 9459 20457
rect 9401 20417 9413 20451
rect 9447 20417 9459 20451
rect 10594 20448 10600 20460
rect 10555 20420 10600 20448
rect 9401 20411 9459 20417
rect 10594 20408 10600 20420
rect 10652 20408 10658 20460
rect 10778 20448 10784 20460
rect 10739 20420 10784 20448
rect 10778 20408 10784 20420
rect 10836 20408 10842 20460
rect 10962 20448 10968 20460
rect 10923 20420 10968 20448
rect 10962 20408 10968 20420
rect 11020 20408 11026 20460
rect 11974 20408 11980 20460
rect 12032 20448 12038 20460
rect 12207 20451 12265 20457
rect 12207 20448 12219 20451
rect 12032 20420 12219 20448
rect 12032 20408 12038 20420
rect 12207 20417 12219 20420
rect 12253 20417 12265 20451
rect 12342 20448 12348 20460
rect 12303 20420 12348 20448
rect 12207 20411 12265 20417
rect 12342 20408 12348 20420
rect 12400 20408 12406 20460
rect 12434 20408 12440 20460
rect 12492 20448 12498 20460
rect 12618 20448 12624 20460
rect 12492 20420 12537 20448
rect 12579 20420 12624 20448
rect 12492 20408 12498 20420
rect 12618 20408 12624 20420
rect 12676 20408 12682 20460
rect 13633 20451 13691 20457
rect 13633 20417 13645 20451
rect 13679 20417 13691 20451
rect 13633 20411 13691 20417
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20417 13783 20451
rect 13725 20411 13783 20417
rect 12066 20340 12072 20392
rect 12124 20380 12130 20392
rect 13648 20380 13676 20411
rect 12124 20352 13676 20380
rect 12124 20340 12130 20352
rect 12250 20312 12256 20324
rect 8404 20284 12256 20312
rect 6362 20204 6368 20256
rect 6420 20244 6426 20256
rect 8404 20244 8432 20284
rect 12250 20272 12256 20284
rect 12308 20272 12314 20324
rect 13740 20312 13768 20411
rect 13814 20408 13820 20460
rect 13872 20448 13878 20460
rect 13872 20420 13917 20448
rect 13872 20408 13878 20420
rect 13998 20408 14004 20460
rect 14056 20448 14062 20460
rect 14752 20457 14780 20488
rect 14737 20451 14795 20457
rect 14056 20420 14101 20448
rect 14056 20408 14062 20420
rect 14737 20417 14749 20451
rect 14783 20417 14795 20451
rect 14737 20411 14795 20417
rect 14826 20451 14884 20457
rect 14826 20417 14838 20451
rect 14872 20417 14884 20451
rect 14826 20411 14884 20417
rect 13906 20312 13912 20324
rect 13740 20284 13912 20312
rect 13906 20272 13912 20284
rect 13964 20312 13970 20324
rect 14844 20312 14872 20411
rect 14918 20408 14924 20460
rect 14976 20448 14982 20460
rect 14976 20420 15021 20448
rect 14976 20408 14982 20420
rect 15102 20408 15108 20460
rect 15160 20448 15166 20460
rect 15657 20451 15715 20457
rect 15160 20420 15205 20448
rect 15160 20408 15166 20420
rect 15657 20417 15669 20451
rect 15703 20417 15715 20451
rect 15657 20411 15715 20417
rect 15672 20380 15700 20411
rect 15838 20408 15844 20460
rect 15896 20448 15902 20460
rect 16758 20448 16764 20460
rect 15896 20420 16764 20448
rect 15896 20408 15902 20420
rect 16758 20408 16764 20420
rect 16816 20408 16822 20460
rect 16940 20457 16968 20488
rect 17678 20476 17684 20488
rect 17736 20476 17742 20528
rect 18233 20519 18291 20525
rect 18233 20485 18245 20519
rect 18279 20516 18291 20519
rect 20254 20516 20260 20528
rect 18279 20488 20260 20516
rect 18279 20485 18291 20488
rect 18233 20479 18291 20485
rect 20254 20476 20260 20488
rect 20312 20476 20318 20528
rect 23768 20516 23796 20556
rect 27982 20516 27988 20528
rect 20548 20488 23796 20516
rect 27943 20488 27988 20516
rect 16940 20451 17003 20457
rect 16940 20420 16957 20451
rect 16945 20417 16957 20420
rect 16991 20417 17003 20451
rect 16945 20411 17003 20417
rect 17037 20451 17095 20457
rect 17037 20417 17049 20451
rect 17083 20417 17095 20451
rect 17037 20411 17095 20417
rect 17129 20451 17187 20457
rect 17129 20417 17141 20451
rect 17175 20417 17187 20451
rect 17129 20411 17187 20417
rect 15930 20380 15936 20392
rect 15672 20352 15936 20380
rect 15930 20340 15936 20352
rect 15988 20340 15994 20392
rect 17052 20312 17080 20411
rect 13964 20284 17080 20312
rect 13964 20272 13970 20284
rect 6420 20216 8432 20244
rect 6420 20204 6426 20216
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11204 20216 11989 20244
rect 11204 20204 11210 20216
rect 11977 20213 11989 20216
rect 12023 20213 12035 20247
rect 11977 20207 12035 20213
rect 13357 20247 13415 20253
rect 13357 20213 13369 20247
rect 13403 20244 13415 20247
rect 13446 20244 13452 20256
rect 13403 20216 13452 20244
rect 13403 20213 13415 20216
rect 13357 20207 13415 20213
rect 13446 20204 13452 20216
rect 13504 20204 13510 20256
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 17144 20244 17172 20411
rect 17310 20408 17316 20460
rect 17368 20448 17374 20460
rect 18046 20448 18052 20460
rect 17368 20420 17413 20448
rect 18007 20420 18052 20448
rect 17368 20408 17374 20420
rect 18046 20408 18052 20420
rect 18104 20408 18110 20460
rect 19613 20451 19671 20457
rect 19613 20417 19625 20451
rect 19659 20448 19671 20451
rect 20070 20448 20076 20460
rect 19659 20420 20076 20448
rect 19659 20417 19671 20420
rect 19613 20411 19671 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20548 20457 20576 20488
rect 27982 20476 27988 20488
rect 28040 20476 28046 20528
rect 28169 20519 28227 20525
rect 28169 20485 28181 20519
rect 28215 20516 28227 20519
rect 29270 20516 29276 20528
rect 28215 20488 29276 20516
rect 28215 20485 28227 20488
rect 28169 20479 28227 20485
rect 29270 20476 29276 20488
rect 29328 20516 29334 20528
rect 29730 20516 29736 20528
rect 29328 20488 29736 20516
rect 29328 20476 29334 20488
rect 29730 20476 29736 20488
rect 29788 20476 29794 20528
rect 31662 20516 31668 20528
rect 30208 20488 31668 20516
rect 30208 20460 30236 20488
rect 31662 20476 31668 20488
rect 31720 20516 31726 20528
rect 34698 20516 34704 20528
rect 31720 20488 34704 20516
rect 31720 20476 31726 20488
rect 20533 20451 20591 20457
rect 20533 20417 20545 20451
rect 20579 20417 20591 20451
rect 20533 20411 20591 20417
rect 20625 20451 20683 20457
rect 20625 20417 20637 20451
rect 20671 20417 20683 20451
rect 20625 20411 20683 20417
rect 18322 20340 18328 20392
rect 18380 20380 18386 20392
rect 19242 20380 19248 20392
rect 18380 20352 19248 20380
rect 18380 20340 18386 20352
rect 19242 20340 19248 20352
rect 19300 20380 19306 20392
rect 20640 20380 20668 20411
rect 20714 20408 20720 20460
rect 20772 20448 20778 20460
rect 20901 20451 20959 20457
rect 20772 20420 20817 20448
rect 20772 20408 20778 20420
rect 20901 20417 20913 20451
rect 20947 20448 20959 20451
rect 20990 20448 20996 20460
rect 20947 20420 20996 20448
rect 20947 20417 20959 20420
rect 20901 20411 20959 20417
rect 20990 20408 20996 20420
rect 21048 20448 21054 20460
rect 22094 20448 22100 20460
rect 21048 20420 22100 20448
rect 21048 20408 21054 20420
rect 22094 20408 22100 20420
rect 22152 20408 22158 20460
rect 23290 20448 23296 20460
rect 23251 20420 23296 20448
rect 23290 20408 23296 20420
rect 23348 20408 23354 20460
rect 23474 20408 23480 20460
rect 23532 20448 23538 20460
rect 30190 20448 30196 20460
rect 23532 20420 28994 20448
rect 30151 20420 30196 20448
rect 23532 20408 23538 20420
rect 19300 20352 20668 20380
rect 19300 20340 19306 20352
rect 21726 20340 21732 20392
rect 21784 20380 21790 20392
rect 23934 20380 23940 20392
rect 21784 20352 23940 20380
rect 21784 20340 21790 20352
rect 23934 20340 23940 20352
rect 23992 20340 23998 20392
rect 17494 20272 17500 20324
rect 17552 20312 17558 20324
rect 26602 20312 26608 20324
rect 17552 20284 26608 20312
rect 17552 20272 17558 20284
rect 26602 20272 26608 20284
rect 26660 20272 26666 20324
rect 17678 20244 17684 20256
rect 16071 20216 17172 20244
rect 17639 20216 17684 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 17678 20204 17684 20216
rect 17736 20204 17742 20256
rect 18417 20247 18475 20253
rect 18417 20213 18429 20247
rect 18463 20244 18475 20247
rect 18506 20244 18512 20256
rect 18463 20216 18512 20244
rect 18463 20213 18475 20216
rect 18417 20207 18475 20213
rect 18506 20204 18512 20216
rect 18564 20204 18570 20256
rect 18598 20204 18604 20256
rect 18656 20244 18662 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 18656 20216 19717 20244
rect 18656 20204 18662 20216
rect 19705 20213 19717 20216
rect 19751 20244 19763 20247
rect 19886 20244 19892 20256
rect 19751 20216 19892 20244
rect 19751 20213 19763 20216
rect 19705 20207 19763 20213
rect 19886 20204 19892 20216
rect 19944 20204 19950 20256
rect 20257 20247 20315 20253
rect 20257 20213 20269 20247
rect 20303 20244 20315 20247
rect 21450 20244 21456 20256
rect 20303 20216 21456 20244
rect 20303 20213 20315 20216
rect 20257 20207 20315 20213
rect 21450 20204 21456 20216
rect 21508 20204 21514 20256
rect 21910 20204 21916 20256
rect 21968 20244 21974 20256
rect 22646 20244 22652 20256
rect 21968 20216 22652 20244
rect 21968 20204 21974 20216
rect 22646 20204 22652 20216
rect 22704 20204 22710 20256
rect 23198 20204 23204 20256
rect 23256 20244 23262 20256
rect 23385 20247 23443 20253
rect 23385 20244 23397 20247
rect 23256 20216 23397 20244
rect 23256 20204 23262 20216
rect 23385 20213 23397 20216
rect 23431 20213 23443 20247
rect 23385 20207 23443 20213
rect 24026 20204 24032 20256
rect 24084 20244 24090 20256
rect 24302 20244 24308 20256
rect 24084 20216 24308 20244
rect 24084 20204 24090 20216
rect 24302 20204 24308 20216
rect 24360 20204 24366 20256
rect 28966 20244 28994 20420
rect 30190 20408 30196 20420
rect 30248 20408 30254 20460
rect 30282 20408 30288 20460
rect 30340 20448 30346 20460
rect 32140 20457 32168 20488
rect 34698 20476 34704 20488
rect 34756 20476 34762 20528
rect 41386 20516 41414 20556
rect 48038 20516 48044 20528
rect 41386 20488 48044 20516
rect 48038 20476 48044 20488
rect 48096 20476 48102 20528
rect 30449 20451 30507 20457
rect 30449 20448 30461 20451
rect 30340 20420 30461 20448
rect 30340 20408 30346 20420
rect 30449 20417 30461 20420
rect 30495 20417 30507 20451
rect 30449 20411 30507 20417
rect 32125 20451 32183 20457
rect 32125 20417 32137 20451
rect 32171 20417 32183 20451
rect 32125 20411 32183 20417
rect 32214 20408 32220 20460
rect 32272 20448 32278 20460
rect 32381 20451 32439 20457
rect 32381 20448 32393 20451
rect 32272 20420 32393 20448
rect 32272 20408 32278 20420
rect 32381 20417 32393 20420
rect 32427 20417 32439 20451
rect 32381 20411 32439 20417
rect 32674 20408 32680 20460
rect 32732 20448 32738 20460
rect 34238 20448 34244 20460
rect 32732 20420 33180 20448
rect 34199 20420 34244 20448
rect 32732 20408 32738 20420
rect 33152 20380 33180 20420
rect 34238 20408 34244 20420
rect 34296 20408 34302 20460
rect 34333 20451 34391 20457
rect 34333 20417 34345 20451
rect 34379 20417 34391 20451
rect 34333 20411 34391 20417
rect 34348 20380 34376 20411
rect 34422 20408 34428 20460
rect 34480 20448 34486 20460
rect 34480 20420 34525 20448
rect 34480 20408 34486 20420
rect 34606 20408 34612 20460
rect 34664 20448 34670 20460
rect 34664 20420 34709 20448
rect 34664 20408 34670 20420
rect 34514 20380 34520 20392
rect 33152 20352 33548 20380
rect 34348 20352 34520 20380
rect 31386 20272 31392 20324
rect 31444 20312 31450 20324
rect 33520 20321 33548 20352
rect 34514 20340 34520 20352
rect 34572 20340 34578 20392
rect 31573 20315 31631 20321
rect 31573 20312 31585 20315
rect 31444 20284 31585 20312
rect 31444 20272 31450 20284
rect 31573 20281 31585 20284
rect 31619 20281 31631 20315
rect 31573 20275 31631 20281
rect 33505 20315 33563 20321
rect 33505 20281 33517 20315
rect 33551 20281 33563 20315
rect 41598 20312 41604 20324
rect 33505 20275 33563 20281
rect 33612 20284 41604 20312
rect 33612 20244 33640 20284
rect 41598 20272 41604 20284
rect 41656 20272 41662 20324
rect 33962 20244 33968 20256
rect 28966 20216 33640 20244
rect 33923 20216 33968 20244
rect 33962 20204 33968 20216
rect 34020 20204 34026 20256
rect 1104 20154 48852 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 48852 20154
rect 1104 20080 48852 20102
rect 10778 20000 10784 20052
rect 10836 20040 10842 20052
rect 11517 20043 11575 20049
rect 11517 20040 11529 20043
rect 10836 20012 11529 20040
rect 10836 20000 10842 20012
rect 11517 20009 11529 20012
rect 11563 20009 11575 20043
rect 11517 20003 11575 20009
rect 13541 20043 13599 20049
rect 13541 20009 13553 20043
rect 13587 20040 13599 20043
rect 13814 20040 13820 20052
rect 13587 20012 13820 20040
rect 13587 20009 13599 20012
rect 13541 20003 13599 20009
rect 13814 20000 13820 20012
rect 13872 20000 13878 20052
rect 14461 20043 14519 20049
rect 14461 20009 14473 20043
rect 14507 20040 14519 20043
rect 14918 20040 14924 20052
rect 14507 20012 14924 20040
rect 14507 20009 14519 20012
rect 14461 20003 14519 20009
rect 14918 20000 14924 20012
rect 14976 20000 14982 20052
rect 15028 20012 17161 20040
rect 12250 19932 12256 19984
rect 12308 19972 12314 19984
rect 15028 19972 15056 20012
rect 12308 19944 15056 19972
rect 17133 19972 17161 20012
rect 17678 20000 17684 20052
rect 17736 20040 17742 20052
rect 47026 20040 47032 20052
rect 17736 20012 47032 20040
rect 17736 20000 17742 20012
rect 47026 20000 47032 20012
rect 47084 20000 47090 20052
rect 17133 19944 18543 19972
rect 12308 19932 12314 19944
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 12342 19904 12348 19916
rect 12124 19876 12348 19904
rect 12124 19864 12130 19876
rect 12342 19864 12348 19876
rect 12400 19904 12406 19916
rect 16114 19904 16120 19916
rect 12400 19876 16120 19904
rect 12400 19864 12406 19876
rect 16114 19864 16120 19876
rect 16172 19904 16178 19916
rect 18515 19904 18543 19944
rect 20254 19932 20260 19984
rect 20312 19972 20318 19984
rect 20530 19972 20536 19984
rect 20312 19944 20536 19972
rect 20312 19932 20318 19944
rect 20530 19932 20536 19944
rect 20588 19972 20594 19984
rect 20625 19975 20683 19981
rect 20625 19972 20637 19975
rect 20588 19944 20637 19972
rect 20588 19932 20594 19944
rect 20625 19941 20637 19944
rect 20671 19941 20683 19975
rect 25774 19972 25780 19984
rect 25735 19944 25780 19972
rect 20625 19935 20683 19941
rect 25774 19932 25780 19944
rect 25832 19932 25838 19984
rect 26513 19975 26571 19981
rect 26513 19941 26525 19975
rect 26559 19972 26571 19975
rect 26786 19972 26792 19984
rect 26559 19944 26792 19972
rect 26559 19941 26571 19944
rect 26513 19935 26571 19941
rect 26786 19932 26792 19944
rect 26844 19932 26850 19984
rect 31202 19932 31208 19984
rect 31260 19972 31266 19984
rect 34057 19975 34115 19981
rect 31260 19944 33916 19972
rect 31260 19932 31266 19944
rect 16172 19876 18460 19904
rect 18515 19876 19380 19904
rect 16172 19864 16178 19876
rect 1854 19796 1860 19848
rect 1912 19836 1918 19848
rect 2041 19839 2099 19845
rect 2041 19836 2053 19839
rect 1912 19808 2053 19836
rect 1912 19796 1918 19808
rect 2041 19805 2053 19808
rect 2087 19805 2099 19839
rect 2041 19799 2099 19805
rect 10137 19839 10195 19845
rect 10137 19805 10149 19839
rect 10183 19805 10195 19839
rect 10137 19799 10195 19805
rect 10404 19839 10462 19845
rect 10404 19805 10416 19839
rect 10450 19836 10462 19839
rect 11146 19836 11152 19848
rect 10450 19808 11152 19836
rect 10450 19805 10462 19808
rect 10404 19799 10462 19805
rect 7834 19728 7840 19780
rect 7892 19768 7898 19780
rect 10152 19768 10180 19799
rect 11146 19796 11152 19808
rect 11204 19796 11210 19848
rect 11790 19796 11796 19848
rect 11848 19836 11854 19848
rect 12161 19839 12219 19845
rect 12161 19836 12173 19839
rect 11848 19808 12173 19836
rect 11848 19796 11854 19808
rect 12161 19805 12173 19808
rect 12207 19805 12219 19839
rect 12161 19799 12219 19805
rect 12986 19796 12992 19848
rect 13044 19836 13050 19848
rect 13173 19839 13231 19845
rect 13173 19836 13185 19839
rect 13044 19808 13185 19836
rect 13044 19796 13050 19808
rect 13173 19805 13185 19808
rect 13219 19836 13231 19839
rect 14274 19836 14280 19848
rect 13219 19808 14136 19836
rect 14235 19808 14280 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 7892 19740 10456 19768
rect 7892 19728 7898 19740
rect 10428 19712 10456 19740
rect 10594 19728 10600 19780
rect 10652 19768 10658 19780
rect 11977 19771 12035 19777
rect 11977 19768 11989 19771
rect 10652 19740 11989 19768
rect 10652 19728 10658 19740
rect 11977 19737 11989 19740
rect 12023 19737 12035 19771
rect 13354 19768 13360 19780
rect 13315 19740 13360 19768
rect 11977 19731 12035 19737
rect 13354 19728 13360 19740
rect 13412 19728 13418 19780
rect 14108 19777 14136 19808
rect 14274 19796 14280 19808
rect 14332 19796 14338 19848
rect 16850 19796 16856 19848
rect 16908 19836 16914 19848
rect 17052 19845 17080 19876
rect 16945 19839 17003 19845
rect 16945 19836 16957 19839
rect 16908 19808 16957 19836
rect 16908 19796 16914 19808
rect 16945 19805 16957 19808
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17037 19839 17095 19845
rect 17037 19805 17049 19839
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 17150 19839 17208 19845
rect 17150 19805 17162 19839
rect 17196 19836 17208 19839
rect 17313 19839 17371 19845
rect 17196 19808 17264 19836
rect 17196 19805 17208 19808
rect 17150 19799 17208 19805
rect 14093 19771 14151 19777
rect 14093 19737 14105 19771
rect 14139 19768 14151 19771
rect 15930 19768 15936 19780
rect 14139 19740 15936 19768
rect 14139 19737 14151 19740
rect 14093 19731 14151 19737
rect 15930 19728 15936 19740
rect 15988 19728 15994 19780
rect 17236 19768 17264 19808
rect 17313 19805 17325 19839
rect 17359 19836 17371 19839
rect 17678 19836 17684 19848
rect 17359 19808 17684 19836
rect 17359 19805 17371 19808
rect 17313 19799 17371 19805
rect 17678 19796 17684 19808
rect 17736 19796 17742 19848
rect 18230 19796 18236 19848
rect 18288 19845 18294 19848
rect 18432 19845 18460 19876
rect 18288 19839 18337 19845
rect 18288 19805 18291 19839
rect 18325 19805 18337 19839
rect 18288 19799 18337 19805
rect 18417 19839 18475 19845
rect 18417 19805 18429 19839
rect 18463 19805 18475 19839
rect 18417 19799 18475 19805
rect 18288 19796 18294 19799
rect 18506 19796 18512 19848
rect 18564 19836 18570 19848
rect 18564 19808 18609 19836
rect 18564 19796 18570 19808
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19242 19836 19248 19848
rect 18748 19808 18793 19836
rect 19203 19808 19248 19836
rect 18748 19796 18754 19808
rect 19242 19796 19248 19808
rect 19300 19796 19306 19848
rect 19352 19836 19380 19876
rect 26602 19864 26608 19916
rect 26660 19904 26666 19916
rect 26660 19876 29684 19904
rect 26660 19864 26666 19876
rect 19352 19808 19656 19836
rect 17494 19768 17500 19780
rect 17236 19740 17500 19768
rect 17494 19728 17500 19740
rect 17552 19728 17558 19780
rect 18049 19771 18107 19777
rect 18049 19737 18061 19771
rect 18095 19737 18107 19771
rect 19490 19771 19548 19777
rect 19490 19768 19502 19771
rect 18049 19731 18107 19737
rect 19306 19740 19502 19768
rect 4062 19660 4068 19712
rect 4120 19700 4126 19712
rect 8202 19700 8208 19712
rect 4120 19672 8208 19700
rect 4120 19660 4126 19672
rect 8202 19660 8208 19672
rect 8260 19660 8266 19712
rect 10410 19660 10416 19712
rect 10468 19660 10474 19712
rect 12345 19703 12403 19709
rect 12345 19669 12357 19703
rect 12391 19700 12403 19703
rect 12802 19700 12808 19712
rect 12391 19672 12808 19700
rect 12391 19669 12403 19672
rect 12345 19663 12403 19669
rect 12802 19660 12808 19672
rect 12860 19660 12866 19712
rect 16669 19703 16727 19709
rect 16669 19669 16681 19703
rect 16715 19700 16727 19703
rect 16850 19700 16856 19712
rect 16715 19672 16856 19700
rect 16715 19669 16727 19672
rect 16669 19663 16727 19669
rect 16850 19660 16856 19672
rect 16908 19660 16914 19712
rect 18064 19700 18092 19731
rect 19306 19700 19334 19740
rect 19490 19737 19502 19740
rect 19536 19737 19548 19771
rect 19628 19768 19656 19808
rect 19886 19796 19892 19848
rect 19944 19836 19950 19848
rect 20254 19836 20260 19848
rect 19944 19808 20260 19836
rect 19944 19796 19950 19808
rect 20254 19796 20260 19808
rect 20312 19796 20318 19848
rect 21174 19836 21180 19848
rect 21135 19808 21180 19836
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21450 19845 21456 19848
rect 21444 19836 21456 19845
rect 21411 19808 21456 19836
rect 21444 19799 21456 19808
rect 21450 19796 21456 19799
rect 21508 19796 21514 19848
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19836 24455 19839
rect 25590 19836 25596 19848
rect 24443 19808 25596 19836
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 25590 19796 25596 19808
rect 25648 19836 25654 19848
rect 27614 19836 27620 19848
rect 25648 19808 27620 19836
rect 25648 19796 25654 19808
rect 27614 19796 27620 19808
rect 27672 19836 27678 19848
rect 27985 19839 28043 19845
rect 27985 19836 27997 19839
rect 27672 19808 27997 19836
rect 27672 19796 27678 19808
rect 27985 19805 27997 19808
rect 28031 19836 28043 19839
rect 29549 19839 29607 19845
rect 29549 19836 29561 19839
rect 28031 19808 29561 19836
rect 28031 19805 28043 19808
rect 27985 19799 28043 19805
rect 29549 19805 29561 19808
rect 29595 19805 29607 19839
rect 29656 19836 29684 19876
rect 31386 19864 31392 19916
rect 31444 19904 31450 19916
rect 31444 19876 31616 19904
rect 31444 19864 31450 19876
rect 30742 19836 30748 19848
rect 29656 19808 30748 19836
rect 29549 19799 29607 19805
rect 30742 19796 30748 19808
rect 30800 19796 30806 19848
rect 31588 19845 31616 19876
rect 33888 19848 33916 19944
rect 34057 19941 34069 19975
rect 34103 19972 34115 19975
rect 34422 19972 34428 19984
rect 34103 19944 34428 19972
rect 34103 19941 34115 19944
rect 34057 19935 34115 19941
rect 34422 19932 34428 19944
rect 34480 19932 34486 19984
rect 34698 19904 34704 19916
rect 34659 19876 34704 19904
rect 34698 19864 34704 19876
rect 34756 19864 34762 19916
rect 46293 19907 46351 19913
rect 46293 19873 46305 19907
rect 46339 19904 46351 19907
rect 47762 19904 47768 19916
rect 46339 19876 47768 19904
rect 46339 19873 46351 19876
rect 46293 19867 46351 19873
rect 47762 19864 47768 19876
rect 47820 19864 47826 19916
rect 31573 19839 31631 19845
rect 31573 19805 31585 19839
rect 31619 19805 31631 19839
rect 32217 19839 32275 19845
rect 32217 19836 32229 19839
rect 31573 19799 31631 19805
rect 31726 19808 32229 19836
rect 24664 19771 24722 19777
rect 19628 19740 24164 19768
rect 19490 19731 19548 19737
rect 22554 19700 22560 19712
rect 18064 19672 19334 19700
rect 22515 19672 22560 19700
rect 22554 19660 22560 19672
rect 22612 19660 22618 19712
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 23658 19700 23664 19712
rect 22704 19672 23664 19700
rect 22704 19660 22710 19672
rect 23658 19660 23664 19672
rect 23716 19660 23722 19712
rect 24136 19700 24164 19740
rect 24664 19737 24676 19771
rect 24710 19768 24722 19771
rect 26050 19768 26056 19780
rect 24710 19740 26056 19768
rect 24710 19737 24722 19740
rect 24664 19731 24722 19737
rect 26050 19728 26056 19740
rect 26108 19728 26114 19780
rect 26329 19771 26387 19777
rect 26329 19737 26341 19771
rect 26375 19737 26387 19771
rect 27798 19768 27804 19780
rect 27759 19740 27804 19768
rect 26329 19731 26387 19737
rect 24762 19700 24768 19712
rect 24136 19672 24768 19700
rect 24762 19660 24768 19672
rect 24820 19700 24826 19712
rect 26344 19700 26372 19731
rect 27798 19728 27804 19740
rect 27856 19728 27862 19780
rect 28626 19728 28632 19780
rect 28684 19768 28690 19780
rect 29794 19771 29852 19777
rect 29794 19768 29806 19771
rect 28684 19740 29806 19768
rect 28684 19728 28690 19740
rect 29794 19737 29806 19740
rect 29840 19737 29852 19771
rect 31389 19771 31447 19777
rect 31389 19768 31401 19771
rect 29794 19731 29852 19737
rect 29932 19740 31401 19768
rect 24820 19672 26372 19700
rect 24820 19660 24826 19672
rect 26786 19660 26792 19712
rect 26844 19700 26850 19712
rect 29932 19700 29960 19740
rect 31389 19737 31401 19740
rect 31435 19768 31447 19771
rect 31726 19768 31754 19808
rect 32217 19805 32229 19808
rect 32263 19836 32275 19839
rect 32306 19836 32312 19848
rect 32263 19808 32312 19836
rect 32263 19805 32275 19808
rect 32217 19799 32275 19805
rect 32306 19796 32312 19808
rect 32364 19796 32370 19848
rect 32401 19839 32459 19845
rect 32401 19805 32413 19839
rect 32447 19836 32459 19839
rect 33226 19836 33232 19848
rect 32447 19808 33232 19836
rect 32447 19805 32459 19808
rect 32401 19799 32459 19805
rect 33226 19796 33232 19808
rect 33284 19796 33290 19848
rect 33686 19836 33692 19848
rect 33647 19808 33692 19836
rect 33686 19796 33692 19808
rect 33744 19796 33750 19848
rect 33870 19836 33876 19848
rect 33783 19808 33876 19836
rect 33870 19796 33876 19808
rect 33928 19796 33934 19848
rect 33962 19796 33968 19848
rect 34020 19836 34026 19848
rect 34957 19839 35015 19845
rect 34957 19836 34969 19839
rect 34020 19808 34969 19836
rect 34020 19796 34026 19808
rect 34957 19805 34969 19808
rect 35003 19805 35015 19839
rect 34957 19799 35015 19805
rect 31435 19740 31754 19768
rect 46477 19771 46535 19777
rect 31435 19737 31447 19740
rect 31389 19731 31447 19737
rect 46477 19737 46489 19771
rect 46523 19768 46535 19771
rect 46750 19768 46756 19780
rect 46523 19740 46756 19768
rect 46523 19737 46535 19740
rect 46477 19731 46535 19737
rect 46750 19728 46756 19740
rect 46808 19728 46814 19780
rect 48130 19768 48136 19780
rect 48091 19740 48136 19768
rect 48130 19728 48136 19740
rect 48188 19728 48194 19780
rect 26844 19672 29960 19700
rect 26844 19660 26850 19672
rect 30006 19660 30012 19712
rect 30064 19700 30070 19712
rect 30929 19703 30987 19709
rect 30929 19700 30941 19703
rect 30064 19672 30941 19700
rect 30064 19660 30070 19672
rect 30929 19669 30941 19672
rect 30975 19669 30987 19703
rect 31754 19700 31760 19712
rect 31715 19672 31760 19700
rect 30929 19663 30987 19669
rect 31754 19660 31760 19672
rect 31812 19660 31818 19712
rect 32030 19660 32036 19712
rect 32088 19700 32094 19712
rect 32585 19703 32643 19709
rect 32585 19700 32597 19703
rect 32088 19672 32597 19700
rect 32088 19660 32094 19672
rect 32585 19669 32597 19672
rect 32631 19669 32643 19703
rect 32585 19663 32643 19669
rect 33870 19660 33876 19712
rect 33928 19700 33934 19712
rect 36081 19703 36139 19709
rect 36081 19700 36093 19703
rect 33928 19672 36093 19700
rect 33928 19660 33934 19672
rect 36081 19669 36093 19672
rect 36127 19669 36139 19703
rect 36081 19663 36139 19669
rect 1104 19610 48852 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 48852 19610
rect 1104 19536 48852 19558
rect 11790 19496 11796 19508
rect 7760 19468 11796 19496
rect 1854 19360 1860 19372
rect 1815 19332 1860 19360
rect 1854 19320 1860 19332
rect 1912 19320 1918 19372
rect 7760 19369 7788 19468
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12434 19456 12440 19508
rect 12492 19456 12498 19508
rect 13354 19456 13360 19508
rect 13412 19496 13418 19508
rect 14553 19499 14611 19505
rect 14553 19496 14565 19499
rect 13412 19468 14565 19496
rect 13412 19456 13418 19468
rect 14553 19465 14565 19468
rect 14599 19465 14611 19499
rect 14553 19459 14611 19465
rect 15102 19456 15108 19508
rect 15160 19496 15166 19508
rect 17310 19496 17316 19508
rect 15160 19468 17316 19496
rect 15160 19456 15166 19468
rect 17310 19456 17316 19468
rect 17368 19456 17374 19508
rect 18138 19496 18144 19508
rect 18051 19468 18144 19496
rect 18138 19456 18144 19468
rect 18196 19496 18202 19508
rect 26050 19496 26056 19508
rect 18196 19468 23060 19496
rect 26011 19468 26056 19496
rect 18196 19456 18202 19468
rect 10781 19431 10839 19437
rect 10781 19397 10793 19431
rect 10827 19428 10839 19431
rect 12158 19428 12164 19440
rect 10827 19400 12164 19428
rect 10827 19397 10839 19400
rect 10781 19391 10839 19397
rect 12158 19388 12164 19400
rect 12216 19388 12222 19440
rect 12452 19375 12480 19456
rect 12802 19428 12808 19440
rect 12636 19400 12808 19428
rect 7745 19363 7803 19369
rect 7745 19329 7757 19363
rect 7791 19329 7803 19363
rect 7745 19323 7803 19329
rect 11974 19320 11980 19372
rect 12032 19360 12038 19372
rect 12450 19369 12508 19375
rect 12345 19363 12403 19369
rect 12345 19360 12357 19363
rect 12032 19332 12357 19360
rect 12032 19320 12038 19332
rect 12345 19329 12357 19332
rect 12391 19329 12403 19363
rect 12450 19335 12462 19369
rect 12496 19335 12508 19369
rect 12450 19329 12508 19335
rect 12550 19363 12608 19369
rect 12550 19329 12562 19363
rect 12596 19360 12608 19363
rect 12636 19360 12664 19400
rect 12802 19388 12808 19400
rect 12860 19388 12866 19440
rect 16114 19428 16120 19440
rect 16075 19400 16120 19428
rect 16114 19388 16120 19400
rect 16172 19388 16178 19440
rect 18877 19431 18935 19437
rect 18877 19428 18889 19431
rect 16776 19400 18889 19428
rect 12596 19332 12664 19360
rect 12596 19329 12608 19332
rect 12345 19323 12403 19329
rect 12550 19323 12608 19329
rect 12710 19320 12716 19372
rect 12768 19360 12774 19372
rect 13170 19360 13176 19372
rect 12768 19332 12813 19360
rect 13131 19332 13176 19360
rect 12768 19320 12793 19332
rect 13170 19320 13176 19332
rect 13228 19320 13234 19372
rect 13446 19369 13452 19372
rect 13440 19360 13452 19369
rect 13407 19332 13452 19360
rect 13440 19323 13452 19332
rect 13446 19320 13452 19323
rect 13504 19320 13510 19372
rect 15838 19320 15844 19372
rect 15896 19360 15902 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15896 19332 15945 19360
rect 15896 19320 15902 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16574 19320 16580 19372
rect 16632 19360 16638 19372
rect 16776 19369 16804 19400
rect 18877 19397 18889 19400
rect 18923 19397 18935 19431
rect 18877 19391 18935 19397
rect 16761 19363 16819 19369
rect 16761 19360 16773 19363
rect 16632 19332 16773 19360
rect 16632 19320 16638 19332
rect 16761 19329 16773 19332
rect 16807 19329 16819 19363
rect 16761 19323 16819 19329
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 17017 19363 17075 19369
rect 17017 19360 17029 19363
rect 16908 19332 17029 19360
rect 16908 19320 16914 19332
rect 17017 19329 17029 19332
rect 17063 19329 17075 19363
rect 17017 19323 17075 19329
rect 17586 19320 17592 19372
rect 17644 19360 17650 19372
rect 18693 19363 18751 19369
rect 18693 19360 18705 19363
rect 17644 19332 18705 19360
rect 17644 19320 17650 19332
rect 18693 19329 18705 19332
rect 18739 19329 18751 19363
rect 18693 19323 18751 19329
rect 12728 19306 12793 19320
rect 2038 19292 2044 19304
rect 1999 19264 2044 19292
rect 2038 19252 2044 19264
rect 2096 19252 2102 19304
rect 2774 19252 2780 19304
rect 2832 19292 2838 19304
rect 7926 19292 7932 19304
rect 2832 19264 2877 19292
rect 7887 19264 7932 19292
rect 2832 19252 2838 19264
rect 7926 19252 7932 19264
rect 7984 19252 7990 19304
rect 8202 19292 8208 19304
rect 8163 19264 8208 19292
rect 8202 19252 8208 19264
rect 8260 19252 8266 19304
rect 10965 19295 11023 19301
rect 10965 19261 10977 19295
rect 11011 19292 11023 19295
rect 12728 19292 12756 19306
rect 11011 19264 12756 19292
rect 18892 19292 18920 19391
rect 19058 19388 19064 19440
rect 19116 19428 19122 19440
rect 19116 19400 20024 19428
rect 19116 19388 19122 19400
rect 19426 19320 19432 19372
rect 19484 19360 19490 19372
rect 19996 19369 20024 19400
rect 20070 19388 20076 19440
rect 20128 19428 20134 19440
rect 22281 19431 22339 19437
rect 22281 19428 22293 19431
rect 20128 19400 22293 19428
rect 20128 19388 20134 19400
rect 22281 19397 22293 19400
rect 22327 19428 22339 19431
rect 22646 19428 22652 19440
rect 22327 19400 22652 19428
rect 22327 19397 22339 19400
rect 22281 19391 22339 19397
rect 22646 19388 22652 19400
rect 22704 19388 22710 19440
rect 19797 19363 19855 19369
rect 19797 19360 19809 19363
rect 19484 19332 19809 19360
rect 19484 19320 19490 19332
rect 19797 19329 19809 19332
rect 19843 19329 19855 19363
rect 19797 19323 19855 19329
rect 19981 19363 20039 19369
rect 19981 19329 19993 19363
rect 20027 19360 20039 19363
rect 22554 19360 22560 19372
rect 20027 19332 22560 19360
rect 20027 19329 20039 19332
rect 19981 19323 20039 19329
rect 22554 19320 22560 19332
rect 22612 19320 22618 19372
rect 23032 19369 23060 19468
rect 26050 19456 26056 19468
rect 26108 19456 26114 19508
rect 28626 19496 28632 19508
rect 28587 19468 28632 19496
rect 28626 19456 28632 19468
rect 28684 19456 28690 19508
rect 30282 19496 30288 19508
rect 30243 19468 30288 19496
rect 30282 19456 30288 19468
rect 30340 19456 30346 19508
rect 30650 19456 30656 19508
rect 30708 19496 30714 19508
rect 31938 19496 31944 19508
rect 30708 19468 31944 19496
rect 30708 19456 30714 19468
rect 31938 19456 31944 19468
rect 31996 19456 32002 19508
rect 32398 19456 32404 19508
rect 32456 19456 32462 19508
rect 33226 19456 33232 19508
rect 33284 19496 33290 19508
rect 33597 19499 33655 19505
rect 33597 19496 33609 19499
rect 33284 19468 33609 19496
rect 33284 19456 33290 19468
rect 33597 19465 33609 19468
rect 33643 19465 33655 19499
rect 46750 19496 46756 19508
rect 46711 19468 46756 19496
rect 33597 19459 33655 19465
rect 46750 19456 46756 19468
rect 46808 19456 46814 19508
rect 23198 19428 23204 19440
rect 23159 19400 23204 19428
rect 23198 19388 23204 19400
rect 23256 19388 23262 19440
rect 23934 19388 23940 19440
rect 23992 19428 23998 19440
rect 23992 19400 29040 19428
rect 23992 19388 23998 19400
rect 23017 19363 23075 19369
rect 23017 19329 23029 19363
rect 23063 19329 23075 19363
rect 23017 19323 23075 19329
rect 25317 19363 25375 19369
rect 25317 19329 25329 19363
rect 25363 19329 25375 19363
rect 25317 19323 25375 19329
rect 21174 19292 21180 19304
rect 18892 19264 21180 19292
rect 11011 19261 11023 19264
rect 10965 19255 11023 19261
rect 21174 19252 21180 19264
rect 21232 19252 21238 19304
rect 23934 19292 23940 19304
rect 23895 19264 23940 19292
rect 23934 19252 23940 19264
rect 23992 19252 23998 19304
rect 24026 19252 24032 19304
rect 24084 19292 24090 19304
rect 25332 19292 25360 19323
rect 25406 19320 25412 19372
rect 25464 19360 25470 19372
rect 26237 19363 26295 19369
rect 26237 19360 26249 19363
rect 25464 19332 26249 19360
rect 25464 19320 25470 19332
rect 26237 19329 26249 19332
rect 26283 19329 26295 19363
rect 28902 19360 28908 19372
rect 28863 19332 28908 19360
rect 26237 19323 26295 19329
rect 28902 19320 28908 19332
rect 28960 19320 28966 19372
rect 29012 19369 29040 19400
rect 30668 19375 30696 19456
rect 31754 19428 31760 19440
rect 30760 19400 31760 19428
rect 28997 19363 29055 19369
rect 28997 19329 29009 19363
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 29086 19320 29092 19372
rect 29144 19360 29150 19372
rect 29144 19332 29189 19360
rect 29144 19320 29150 19332
rect 29270 19320 29276 19372
rect 29328 19360 29334 19372
rect 29328 19332 29373 19360
rect 29328 19320 29334 19332
rect 30006 19320 30012 19372
rect 30064 19360 30070 19372
rect 30650 19369 30708 19375
rect 30760 19369 30788 19400
rect 31754 19388 31760 19400
rect 31812 19388 31818 19440
rect 32416 19428 32444 19456
rect 32416 19400 41414 19428
rect 30515 19363 30573 19369
rect 30515 19360 30527 19363
rect 30064 19332 30527 19360
rect 30064 19320 30070 19332
rect 30515 19329 30527 19332
rect 30561 19329 30573 19363
rect 30650 19335 30662 19369
rect 30696 19335 30708 19369
rect 30650 19329 30708 19335
rect 30745 19363 30803 19369
rect 30745 19329 30757 19363
rect 30791 19329 30803 19363
rect 30515 19323 30573 19329
rect 30745 19323 30803 19329
rect 30929 19363 30987 19369
rect 30929 19329 30941 19363
rect 30975 19360 30987 19363
rect 30975 19332 31616 19360
rect 30975 19329 30987 19332
rect 30929 19323 30987 19329
rect 24084 19264 25360 19292
rect 25593 19295 25651 19301
rect 24084 19252 24090 19264
rect 25593 19261 25605 19295
rect 25639 19292 25651 19295
rect 26418 19292 26424 19304
rect 25639 19264 26424 19292
rect 25639 19261 25651 19264
rect 25593 19255 25651 19261
rect 26418 19252 26424 19264
rect 26476 19252 26482 19304
rect 31588 19292 31616 19332
rect 31662 19320 31668 19372
rect 31720 19360 31726 19372
rect 32217 19363 32275 19369
rect 32217 19360 32229 19363
rect 31720 19332 32229 19360
rect 31720 19320 31726 19332
rect 32217 19329 32229 19332
rect 32263 19329 32275 19363
rect 32217 19323 32275 19329
rect 32306 19320 32312 19372
rect 32364 19360 32370 19372
rect 32473 19363 32531 19369
rect 32473 19360 32485 19363
rect 32364 19332 32485 19360
rect 32364 19320 32370 19332
rect 32473 19329 32485 19332
rect 32519 19329 32531 19363
rect 41386 19360 41414 19400
rect 46661 19363 46719 19369
rect 46661 19360 46673 19363
rect 41386 19332 46673 19360
rect 32473 19323 32531 19329
rect 46661 19329 46673 19332
rect 46707 19329 46719 19363
rect 46661 19323 46719 19329
rect 47762 19292 47768 19304
rect 31588 19264 31754 19292
rect 47723 19264 47768 19292
rect 3510 19184 3516 19236
rect 3568 19224 3574 19236
rect 12894 19224 12900 19236
rect 3568 19196 12900 19224
rect 3568 19184 3574 19196
rect 12894 19184 12900 19196
rect 12952 19184 12958 19236
rect 20165 19227 20223 19233
rect 20165 19193 20177 19227
rect 20211 19224 20223 19227
rect 20714 19224 20720 19236
rect 20211 19196 20720 19224
rect 20211 19193 20223 19196
rect 20165 19187 20223 19193
rect 20714 19184 20720 19196
rect 20772 19184 20778 19236
rect 28626 19224 28632 19236
rect 22388 19196 28632 19224
rect 12066 19156 12072 19168
rect 12027 19128 12072 19156
rect 12066 19116 12072 19128
rect 12124 19116 12130 19168
rect 20530 19116 20536 19168
rect 20588 19156 20594 19168
rect 22186 19156 22192 19168
rect 20588 19128 22192 19156
rect 20588 19116 20594 19128
rect 22186 19116 22192 19128
rect 22244 19116 22250 19168
rect 22278 19116 22284 19168
rect 22336 19156 22342 19168
rect 22388 19165 22416 19196
rect 28626 19184 28632 19196
rect 28684 19184 28690 19236
rect 31726 19224 31754 19264
rect 47762 19252 47768 19264
rect 47820 19252 47826 19304
rect 32214 19224 32220 19236
rect 31726 19196 32220 19224
rect 32214 19184 32220 19196
rect 32272 19184 32278 19236
rect 22373 19159 22431 19165
rect 22373 19156 22385 19159
rect 22336 19128 22385 19156
rect 22336 19116 22342 19128
rect 22373 19125 22385 19128
rect 22419 19125 22431 19159
rect 22373 19119 22431 19125
rect 24670 19116 24676 19168
rect 24728 19156 24734 19168
rect 25409 19159 25467 19165
rect 25409 19156 25421 19159
rect 24728 19128 25421 19156
rect 24728 19116 24734 19128
rect 25409 19125 25421 19128
rect 25455 19125 25467 19159
rect 25409 19119 25467 19125
rect 25501 19159 25559 19165
rect 25501 19125 25513 19159
rect 25547 19156 25559 19159
rect 26602 19156 26608 19168
rect 25547 19128 26608 19156
rect 25547 19125 25559 19128
rect 25501 19119 25559 19125
rect 26602 19116 26608 19128
rect 26660 19116 26666 19168
rect 1104 19066 48852 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 48852 19066
rect 1104 18992 48852 19014
rect 2038 18912 2044 18964
rect 2096 18952 2102 18964
rect 2317 18955 2375 18961
rect 2317 18952 2329 18955
rect 2096 18924 2329 18952
rect 2096 18912 2102 18924
rect 2317 18921 2329 18924
rect 2363 18921 2375 18955
rect 2317 18915 2375 18921
rect 7926 18912 7932 18964
rect 7984 18952 7990 18964
rect 8113 18955 8171 18961
rect 8113 18952 8125 18955
rect 7984 18924 8125 18952
rect 7984 18912 7990 18924
rect 8113 18921 8125 18924
rect 8159 18921 8171 18955
rect 8113 18915 8171 18921
rect 9306 18912 9312 18964
rect 9364 18952 9370 18964
rect 11790 18952 11796 18964
rect 9364 18924 11376 18952
rect 11751 18924 11796 18952
rect 9364 18912 9370 18924
rect 9398 18844 9404 18896
rect 9456 18884 9462 18896
rect 9456 18856 9628 18884
rect 9456 18844 9462 18856
rect 3786 18816 3792 18828
rect 2746 18788 3792 18816
rect 2225 18751 2283 18757
rect 2225 18717 2237 18751
rect 2271 18748 2283 18751
rect 2746 18748 2774 18788
rect 3786 18776 3792 18788
rect 3844 18816 3850 18828
rect 7742 18816 7748 18828
rect 3844 18788 7748 18816
rect 3844 18776 3850 18788
rect 7742 18776 7748 18788
rect 7800 18776 7806 18828
rect 8294 18776 8300 18828
rect 8352 18816 8358 18828
rect 8352 18788 9444 18816
rect 8352 18776 8358 18788
rect 7098 18748 7104 18760
rect 2271 18720 2774 18748
rect 7059 18720 7104 18748
rect 2271 18717 2283 18720
rect 2225 18711 2283 18717
rect 7098 18708 7104 18720
rect 7156 18708 7162 18760
rect 8018 18748 8024 18760
rect 7931 18720 8024 18748
rect 8018 18708 8024 18720
rect 8076 18708 8082 18760
rect 8662 18708 8668 18760
rect 8720 18748 8726 18760
rect 9416 18757 9444 18788
rect 9600 18760 9628 18856
rect 9217 18751 9275 18757
rect 9217 18748 9229 18751
rect 8720 18720 9229 18748
rect 8720 18708 8726 18720
rect 9217 18717 9229 18720
rect 9263 18717 9275 18751
rect 9217 18711 9275 18717
rect 9309 18751 9367 18757
rect 9309 18717 9321 18751
rect 9355 18717 9367 18751
rect 9309 18711 9367 18717
rect 9401 18751 9459 18757
rect 9401 18717 9413 18751
rect 9447 18717 9459 18751
rect 9401 18711 9459 18717
rect 8036 18680 8064 18708
rect 9324 18680 9352 18711
rect 9582 18708 9588 18760
rect 9640 18748 9646 18760
rect 9640 18720 9685 18748
rect 9640 18708 9646 18720
rect 9968 18680 9996 18924
rect 11348 18884 11376 18924
rect 11790 18912 11796 18924
rect 11848 18912 11854 18964
rect 11974 18912 11980 18964
rect 12032 18952 12038 18964
rect 13354 18952 13360 18964
rect 12032 18924 13360 18952
rect 12032 18912 12038 18924
rect 13354 18912 13360 18924
rect 13412 18912 13418 18964
rect 17494 18912 17500 18964
rect 17552 18952 17558 18964
rect 17589 18955 17647 18961
rect 17589 18952 17601 18955
rect 17552 18924 17601 18952
rect 17552 18912 17558 18924
rect 17589 18921 17601 18924
rect 17635 18921 17647 18955
rect 17589 18915 17647 18921
rect 24765 18955 24823 18961
rect 24765 18921 24777 18955
rect 24811 18952 24823 18955
rect 25406 18952 25412 18964
rect 24811 18924 25412 18952
rect 24811 18921 24823 18924
rect 24765 18915 24823 18921
rect 25406 18912 25412 18924
rect 25464 18912 25470 18964
rect 26418 18952 26424 18964
rect 26379 18924 26424 18952
rect 26418 18912 26424 18924
rect 26476 18912 26482 18964
rect 28997 18955 29055 18961
rect 28997 18921 29009 18955
rect 29043 18952 29055 18955
rect 29086 18952 29092 18964
rect 29043 18924 29092 18952
rect 29043 18921 29055 18924
rect 28997 18915 29055 18921
rect 29086 18912 29092 18924
rect 29144 18912 29150 18964
rect 30101 18955 30159 18961
rect 30101 18921 30113 18955
rect 30147 18952 30159 18955
rect 30190 18952 30196 18964
rect 30147 18924 30196 18952
rect 30147 18921 30159 18924
rect 30101 18915 30159 18921
rect 30190 18912 30196 18924
rect 30248 18912 30254 18964
rect 31573 18955 31631 18961
rect 31573 18921 31585 18955
rect 31619 18952 31631 18955
rect 32306 18952 32312 18964
rect 31619 18924 32312 18952
rect 31619 18921 31631 18924
rect 31573 18915 31631 18921
rect 32306 18912 32312 18924
rect 32364 18912 32370 18964
rect 15654 18884 15660 18896
rect 11348 18856 15660 18884
rect 15654 18844 15660 18856
rect 15712 18844 15718 18896
rect 25866 18844 25872 18896
rect 25924 18884 25930 18896
rect 26234 18884 26240 18896
rect 25924 18856 26240 18884
rect 25924 18844 25930 18856
rect 26234 18844 26240 18856
rect 26292 18884 26298 18896
rect 26292 18856 26556 18884
rect 26292 18844 26298 18856
rect 12250 18816 12256 18828
rect 12211 18788 12256 18816
rect 12250 18776 12256 18788
rect 12308 18776 12314 18828
rect 18046 18816 18052 18828
rect 17236 18788 18052 18816
rect 10410 18748 10416 18760
rect 10371 18720 10416 18748
rect 10410 18708 10416 18720
rect 10468 18708 10474 18760
rect 10680 18751 10738 18757
rect 10680 18717 10692 18751
rect 10726 18748 10738 18751
rect 12066 18748 12072 18760
rect 10726 18720 12072 18748
rect 10726 18717 10738 18720
rect 10680 18711 10738 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12434 18708 12440 18760
rect 12492 18748 12498 18760
rect 12529 18751 12587 18757
rect 12529 18748 12541 18751
rect 12492 18720 12541 18748
rect 12492 18708 12498 18720
rect 12529 18717 12541 18720
rect 12575 18717 12587 18751
rect 15746 18748 15752 18760
rect 15707 18720 15752 18748
rect 12529 18711 12587 18717
rect 15746 18708 15752 18720
rect 15804 18708 15810 18760
rect 17236 18757 17264 18788
rect 18046 18776 18052 18788
rect 18104 18776 18110 18828
rect 22646 18776 22652 18828
rect 22704 18816 22710 18828
rect 22741 18819 22799 18825
rect 22741 18816 22753 18819
rect 22704 18788 22753 18816
rect 22704 18776 22710 18788
rect 22741 18785 22753 18788
rect 22787 18785 22799 18819
rect 22741 18779 22799 18785
rect 25317 18819 25375 18825
rect 25317 18785 25329 18819
rect 25363 18816 25375 18819
rect 25363 18788 25544 18816
rect 25363 18785 25375 18788
rect 25317 18779 25375 18785
rect 16025 18751 16083 18757
rect 16025 18717 16037 18751
rect 16071 18748 16083 18751
rect 17221 18751 17279 18757
rect 17221 18748 17233 18751
rect 16071 18720 17233 18748
rect 16071 18717 16083 18720
rect 16025 18711 16083 18717
rect 17221 18717 17233 18720
rect 17267 18717 17279 18751
rect 17221 18711 17279 18717
rect 17405 18751 17463 18757
rect 17405 18717 17417 18751
rect 17451 18748 17463 18751
rect 18138 18748 18144 18760
rect 17451 18720 18144 18748
rect 17451 18717 17463 18720
rect 17405 18711 17463 18717
rect 8036 18652 9076 18680
rect 9324 18652 9996 18680
rect 6822 18572 6828 18624
rect 6880 18612 6886 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 6880 18584 7205 18612
rect 6880 18572 6886 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 8938 18612 8944 18624
rect 8899 18584 8944 18612
rect 7193 18575 7251 18581
rect 8938 18572 8944 18584
rect 8996 18572 9002 18624
rect 9048 18612 9076 18652
rect 10594 18640 10600 18692
rect 10652 18680 10658 18692
rect 16040 18680 16068 18711
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 22462 18748 22468 18760
rect 22423 18720 22468 18748
rect 22462 18708 22468 18720
rect 22520 18708 22526 18760
rect 22557 18751 22615 18757
rect 22557 18717 22569 18751
rect 22603 18748 22615 18751
rect 24670 18748 24676 18760
rect 22603 18720 24676 18748
rect 22603 18717 22615 18720
rect 22557 18711 22615 18717
rect 24670 18708 24676 18720
rect 24728 18708 24734 18760
rect 24946 18708 24952 18760
rect 25004 18748 25010 18760
rect 25406 18748 25412 18760
rect 25004 18720 25412 18748
rect 25004 18708 25010 18720
rect 25406 18708 25412 18720
rect 25464 18708 25470 18760
rect 25516 18748 25544 18788
rect 26142 18748 26148 18760
rect 25516 18720 25912 18748
rect 26103 18720 26148 18748
rect 25130 18680 25136 18692
rect 10652 18652 16068 18680
rect 25043 18652 25136 18680
rect 10652 18640 10658 18652
rect 25130 18640 25136 18652
rect 25188 18680 25194 18692
rect 25774 18680 25780 18692
rect 25188 18652 25780 18680
rect 25188 18640 25194 18652
rect 25774 18640 25780 18652
rect 25832 18640 25838 18692
rect 25884 18680 25912 18720
rect 26142 18708 26148 18720
rect 26200 18708 26206 18760
rect 26528 18757 26556 18856
rect 28902 18844 28908 18896
rect 28960 18884 28966 18896
rect 28960 18856 47624 18884
rect 28960 18844 28966 18856
rect 28718 18776 28724 18828
rect 28776 18816 28782 18828
rect 47302 18816 47308 18828
rect 28776 18788 41414 18816
rect 47263 18788 47308 18816
rect 28776 18776 28782 18788
rect 26237 18751 26295 18757
rect 26237 18717 26249 18751
rect 26283 18717 26295 18751
rect 26237 18711 26295 18717
rect 26513 18751 26571 18757
rect 26513 18717 26525 18751
rect 26559 18717 26571 18751
rect 26513 18711 26571 18717
rect 26252 18680 26280 18711
rect 27798 18708 27804 18760
rect 27856 18748 27862 18760
rect 28169 18751 28227 18757
rect 28169 18748 28181 18751
rect 27856 18720 28181 18748
rect 27856 18708 27862 18720
rect 28169 18717 28181 18720
rect 28215 18748 28227 18751
rect 30009 18751 30067 18757
rect 30009 18748 30021 18751
rect 28215 18720 30021 18748
rect 28215 18717 28227 18720
rect 28169 18711 28227 18717
rect 30009 18717 30021 18720
rect 30055 18717 30067 18751
rect 31846 18748 31852 18760
rect 31807 18720 31852 18748
rect 30009 18711 30067 18717
rect 31846 18708 31852 18720
rect 31904 18708 31910 18760
rect 31941 18751 31999 18757
rect 31941 18717 31953 18751
rect 31987 18717 31999 18751
rect 31941 18711 31999 18717
rect 26602 18680 26608 18692
rect 25884 18652 26096 18680
rect 26252 18652 26608 18680
rect 11882 18612 11888 18624
rect 9048 18584 11888 18612
rect 11882 18572 11888 18584
rect 11940 18572 11946 18624
rect 22741 18615 22799 18621
rect 22741 18581 22753 18615
rect 22787 18612 22799 18615
rect 23658 18612 23664 18624
rect 22787 18584 23664 18612
rect 22787 18581 22799 18584
rect 22741 18575 22799 18581
rect 23658 18572 23664 18584
rect 23716 18572 23722 18624
rect 24394 18572 24400 18624
rect 24452 18612 24458 18624
rect 24578 18612 24584 18624
rect 24452 18584 24584 18612
rect 24452 18572 24458 18584
rect 24578 18572 24584 18584
rect 24636 18572 24642 18624
rect 25225 18615 25283 18621
rect 25225 18581 25237 18615
rect 25271 18612 25283 18615
rect 25961 18615 26019 18621
rect 25961 18612 25973 18615
rect 25271 18584 25973 18612
rect 25271 18581 25283 18584
rect 25225 18575 25283 18581
rect 25961 18581 25973 18584
rect 26007 18581 26019 18615
rect 26068 18612 26096 18652
rect 26602 18640 26608 18652
rect 26660 18640 26666 18692
rect 27982 18680 27988 18692
rect 27943 18652 27988 18680
rect 27982 18640 27988 18652
rect 28040 18640 28046 18692
rect 28626 18680 28632 18692
rect 28587 18652 28632 18680
rect 28626 18640 28632 18652
rect 28684 18640 28690 18692
rect 28813 18683 28871 18689
rect 28813 18649 28825 18683
rect 28859 18680 28871 18683
rect 29914 18680 29920 18692
rect 28859 18652 29920 18680
rect 28859 18649 28871 18652
rect 28813 18643 28871 18649
rect 29914 18640 29920 18652
rect 29972 18640 29978 18692
rect 31956 18624 31984 18711
rect 32030 18708 32036 18760
rect 32088 18748 32094 18760
rect 32088 18720 32133 18748
rect 32088 18708 32094 18720
rect 32214 18708 32220 18760
rect 32272 18748 32278 18760
rect 32582 18748 32588 18760
rect 32272 18720 32588 18748
rect 32272 18708 32278 18720
rect 32582 18708 32588 18720
rect 32640 18708 32646 18760
rect 41386 18748 41414 18788
rect 47302 18776 47308 18788
rect 47360 18776 47366 18828
rect 47596 18825 47624 18856
rect 47581 18819 47639 18825
rect 47581 18785 47593 18819
rect 47627 18785 47639 18819
rect 47581 18779 47639 18785
rect 46198 18748 46204 18760
rect 41386 18720 46204 18748
rect 46198 18708 46204 18720
rect 46256 18708 46262 18760
rect 29270 18612 29276 18624
rect 26068 18584 29276 18612
rect 25961 18575 26019 18581
rect 29270 18572 29276 18584
rect 29328 18572 29334 18624
rect 31938 18572 31944 18624
rect 31996 18572 32002 18624
rect 1104 18522 48852 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 48852 18522
rect 1104 18448 48852 18470
rect 7834 18408 7840 18420
rect 6748 18380 7840 18408
rect 6748 18349 6776 18380
rect 7834 18368 7840 18380
rect 7892 18368 7898 18420
rect 22094 18408 22100 18420
rect 7944 18380 22100 18408
rect 6733 18343 6791 18349
rect 6733 18309 6745 18343
rect 6779 18309 6791 18343
rect 6733 18303 6791 18309
rect 6822 18300 6828 18352
rect 6880 18340 6886 18352
rect 6880 18312 6925 18340
rect 6880 18300 6886 18312
rect 2041 18275 2099 18281
rect 2041 18241 2053 18275
rect 2087 18241 2099 18275
rect 2682 18272 2688 18284
rect 2643 18244 2688 18272
rect 2041 18235 2099 18241
rect 2056 18204 2084 18235
rect 2682 18232 2688 18244
rect 2740 18232 2746 18284
rect 7944 18272 7972 18380
rect 22094 18368 22100 18380
rect 22152 18368 22158 18420
rect 24670 18368 24676 18420
rect 24728 18408 24734 18420
rect 25133 18411 25191 18417
rect 25133 18408 25145 18411
rect 24728 18380 25145 18408
rect 24728 18368 24734 18380
rect 25133 18377 25145 18380
rect 25179 18377 25191 18411
rect 25133 18371 25191 18377
rect 25593 18411 25651 18417
rect 25593 18377 25605 18411
rect 25639 18377 25651 18411
rect 25593 18371 25651 18377
rect 8104 18343 8162 18349
rect 8104 18309 8116 18343
rect 8150 18340 8162 18343
rect 8938 18340 8944 18352
rect 8150 18312 8944 18340
rect 8150 18309 8162 18312
rect 8104 18303 8162 18309
rect 8938 18300 8944 18312
rect 8996 18300 9002 18352
rect 10594 18340 10600 18352
rect 10555 18312 10600 18340
rect 10594 18300 10600 18312
rect 10652 18300 10658 18352
rect 10962 18340 10968 18352
rect 10923 18312 10968 18340
rect 10962 18300 10968 18312
rect 11020 18300 11026 18352
rect 15102 18340 15108 18352
rect 14108 18312 15108 18340
rect 7576 18244 7972 18272
rect 10781 18275 10839 18281
rect 2314 18204 2320 18216
rect 2056 18176 2320 18204
rect 2314 18164 2320 18176
rect 2372 18204 2378 18216
rect 7576 18204 7604 18244
rect 10781 18241 10793 18275
rect 10827 18272 10839 18275
rect 10870 18272 10876 18284
rect 10827 18244 10876 18272
rect 10827 18241 10839 18244
rect 10781 18235 10839 18241
rect 10870 18232 10876 18244
rect 10928 18232 10934 18284
rect 11974 18232 11980 18284
rect 12032 18281 12038 18284
rect 12032 18275 12081 18281
rect 12032 18241 12035 18275
rect 12069 18241 12081 18275
rect 12032 18235 12081 18241
rect 12158 18278 12216 18284
rect 12158 18244 12170 18278
rect 12204 18244 12216 18278
rect 12158 18238 12216 18244
rect 12032 18232 12038 18235
rect 7834 18204 7840 18216
rect 2372 18176 7604 18204
rect 7795 18176 7840 18204
rect 2372 18164 2378 18176
rect 7834 18164 7840 18176
rect 7892 18164 7898 18216
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12176 18204 12204 18238
rect 12250 18232 12256 18284
rect 12308 18275 12314 18284
rect 12308 18247 12350 18275
rect 12434 18272 12440 18284
rect 12308 18232 12314 18247
rect 12406 18232 12440 18272
rect 12492 18272 12498 18284
rect 12492 18244 12537 18272
rect 12492 18232 12498 18244
rect 12894 18232 12900 18284
rect 12952 18272 12958 18284
rect 14108 18281 14136 18312
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 15654 18340 15660 18352
rect 15615 18312 15660 18340
rect 15654 18300 15660 18312
rect 15712 18300 15718 18352
rect 16761 18343 16819 18349
rect 16761 18309 16773 18343
rect 16807 18340 16819 18343
rect 17586 18340 17592 18352
rect 16807 18312 17592 18340
rect 16807 18309 16819 18312
rect 16761 18303 16819 18309
rect 17586 18300 17592 18312
rect 17644 18300 17650 18352
rect 19153 18343 19211 18349
rect 19153 18309 19165 18343
rect 19199 18340 19211 18343
rect 19426 18340 19432 18352
rect 19199 18312 19432 18340
rect 19199 18309 19211 18312
rect 19153 18303 19211 18309
rect 19426 18300 19432 18312
rect 19484 18300 19490 18352
rect 25608 18340 25636 18371
rect 25774 18368 25780 18420
rect 25832 18408 25838 18420
rect 26053 18411 26111 18417
rect 26053 18408 26065 18411
rect 25832 18380 26065 18408
rect 25832 18368 25838 18380
rect 26053 18377 26065 18380
rect 26099 18377 26111 18411
rect 26053 18371 26111 18377
rect 25866 18340 25872 18352
rect 24780 18312 25872 18340
rect 13679 18275 13737 18281
rect 13679 18272 13691 18275
rect 12952 18244 13691 18272
rect 12952 18232 12958 18244
rect 13679 18241 13691 18244
rect 13725 18241 13737 18275
rect 13679 18235 13737 18241
rect 13830 18275 13888 18281
rect 13830 18241 13842 18275
rect 13876 18241 13888 18275
rect 13830 18235 13888 18241
rect 13930 18275 13988 18281
rect 13930 18241 13942 18275
rect 13976 18272 13988 18275
rect 14093 18275 14151 18281
rect 13976 18244 14044 18272
rect 13976 18241 13988 18244
rect 13930 18235 13988 18241
rect 11848 18176 12204 18204
rect 11848 18164 11854 18176
rect 3142 18096 3148 18148
rect 3200 18136 3206 18148
rect 7285 18139 7343 18145
rect 7285 18136 7297 18139
rect 3200 18108 7297 18136
rect 3200 18096 3206 18108
rect 7285 18105 7297 18108
rect 7331 18105 7343 18139
rect 7285 18099 7343 18105
rect 9582 18096 9588 18148
rect 9640 18136 9646 18148
rect 12406 18136 12434 18232
rect 13845 18204 13873 18235
rect 13845 18176 13952 18204
rect 13924 18148 13952 18176
rect 14016 18148 14044 18244
rect 14093 18241 14105 18275
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14182 18232 14188 18284
rect 14240 18272 14246 18284
rect 14550 18272 14556 18284
rect 14240 18244 14556 18272
rect 14240 18232 14246 18244
rect 14550 18232 14556 18244
rect 14608 18272 14614 18284
rect 14645 18275 14703 18281
rect 14645 18272 14657 18275
rect 14608 18244 14657 18272
rect 14608 18232 14614 18244
rect 14645 18241 14657 18244
rect 14691 18241 14703 18275
rect 14645 18235 14703 18241
rect 15473 18275 15531 18281
rect 15473 18241 15485 18275
rect 15519 18272 15531 18275
rect 15838 18272 15844 18284
rect 15519 18244 15844 18272
rect 15519 18241 15531 18244
rect 15473 18235 15531 18241
rect 15838 18232 15844 18244
rect 15896 18232 15902 18284
rect 17954 18232 17960 18284
rect 18012 18272 18018 18284
rect 18233 18278 18291 18281
rect 18156 18275 18291 18278
rect 18156 18272 18245 18275
rect 18012 18250 18245 18272
rect 18012 18244 18184 18250
rect 18012 18232 18018 18244
rect 18233 18241 18245 18250
rect 18279 18241 18291 18275
rect 18233 18235 18291 18241
rect 18322 18275 18380 18281
rect 18322 18241 18334 18275
rect 18368 18241 18380 18275
rect 18322 18235 18380 18241
rect 18438 18275 18496 18281
rect 18438 18241 18450 18275
rect 18484 18272 18496 18275
rect 18601 18275 18659 18281
rect 18484 18244 18552 18272
rect 18484 18241 18496 18244
rect 18438 18235 18496 18241
rect 18340 18204 18368 18235
rect 18340 18176 18460 18204
rect 18432 18148 18460 18176
rect 9640 18108 12434 18136
rect 9640 18096 9646 18108
rect 13262 18096 13268 18148
rect 13320 18136 13326 18148
rect 13320 18108 13860 18136
rect 13320 18096 13326 18108
rect 1578 18068 1584 18080
rect 1539 18040 1584 18068
rect 1578 18028 1584 18040
rect 1636 18028 1642 18080
rect 2130 18068 2136 18080
rect 2091 18040 2136 18068
rect 2130 18028 2136 18040
rect 2188 18028 2194 18080
rect 2777 18071 2835 18077
rect 2777 18037 2789 18071
rect 2823 18068 2835 18071
rect 2866 18068 2872 18080
rect 2823 18040 2872 18068
rect 2823 18037 2835 18040
rect 2777 18031 2835 18037
rect 2866 18028 2872 18040
rect 2924 18028 2930 18080
rect 8754 18028 8760 18080
rect 8812 18068 8818 18080
rect 9217 18071 9275 18077
rect 9217 18068 9229 18071
rect 8812 18040 9229 18068
rect 8812 18028 8818 18040
rect 9217 18037 9229 18040
rect 9263 18037 9275 18071
rect 11790 18068 11796 18080
rect 11751 18040 11796 18068
rect 9217 18031 9275 18037
rect 11790 18028 11796 18040
rect 11848 18028 11854 18080
rect 11882 18028 11888 18080
rect 11940 18068 11946 18080
rect 12894 18068 12900 18080
rect 11940 18040 12900 18068
rect 11940 18028 11946 18040
rect 12894 18028 12900 18040
rect 12952 18028 12958 18080
rect 13446 18068 13452 18080
rect 13407 18040 13452 18068
rect 13446 18028 13452 18040
rect 13504 18028 13510 18080
rect 13832 18068 13860 18108
rect 13906 18096 13912 18148
rect 13964 18096 13970 18148
rect 13998 18096 14004 18148
rect 14056 18096 14062 18148
rect 18414 18096 18420 18148
rect 18472 18096 18478 18148
rect 18524 18136 18552 18244
rect 18601 18241 18613 18275
rect 18647 18272 18659 18275
rect 18782 18272 18788 18284
rect 18647 18244 18788 18272
rect 18647 18241 18659 18244
rect 18601 18235 18659 18241
rect 18782 18232 18788 18244
rect 18840 18232 18846 18284
rect 19337 18275 19395 18281
rect 19337 18241 19349 18275
rect 19383 18272 19395 18275
rect 20622 18272 20628 18284
rect 19383 18244 20628 18272
rect 19383 18241 19395 18244
rect 19337 18235 19395 18241
rect 20622 18232 20628 18244
rect 20680 18232 20686 18284
rect 21174 18232 21180 18284
rect 21232 18272 21238 18284
rect 21821 18275 21879 18281
rect 21821 18272 21833 18275
rect 21232 18244 21833 18272
rect 21232 18232 21238 18244
rect 21821 18241 21833 18244
rect 21867 18241 21879 18275
rect 21821 18235 21879 18241
rect 22088 18275 22146 18281
rect 22088 18241 22100 18275
rect 22134 18272 22146 18275
rect 23198 18272 23204 18284
rect 22134 18244 23204 18272
rect 22134 18241 22146 18244
rect 22088 18235 22146 18241
rect 23198 18232 23204 18244
rect 23256 18232 23262 18284
rect 23474 18232 23480 18284
rect 23532 18272 23538 18284
rect 24780 18281 24808 18312
rect 25866 18300 25872 18312
rect 25924 18300 25930 18352
rect 23661 18275 23719 18281
rect 23661 18272 23673 18275
rect 23532 18244 23673 18272
rect 23532 18232 23538 18244
rect 23661 18241 23673 18244
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 24765 18275 24823 18281
rect 24765 18241 24777 18275
rect 24811 18241 24823 18275
rect 24946 18272 24952 18284
rect 24907 18244 24952 18272
rect 24765 18235 24823 18241
rect 24946 18232 24952 18244
rect 25004 18232 25010 18284
rect 25314 18232 25320 18284
rect 25372 18272 25378 18284
rect 25961 18275 26019 18281
rect 25961 18272 25973 18275
rect 25372 18244 25973 18272
rect 25372 18232 25378 18244
rect 25961 18241 25973 18244
rect 26007 18272 26019 18275
rect 26234 18272 26240 18284
rect 26007 18244 26240 18272
rect 26007 18241 26019 18244
rect 25961 18235 26019 18241
rect 26234 18232 26240 18244
rect 26292 18232 26298 18284
rect 27614 18272 27620 18284
rect 27575 18244 27620 18272
rect 27614 18232 27620 18244
rect 27672 18232 27678 18284
rect 27884 18275 27942 18281
rect 27884 18241 27896 18275
rect 27930 18272 27942 18275
rect 28258 18272 28264 18284
rect 27930 18244 28264 18272
rect 27930 18241 27942 18244
rect 27884 18235 27942 18241
rect 28258 18232 28264 18244
rect 28316 18232 28322 18284
rect 23753 18207 23811 18213
rect 23753 18173 23765 18207
rect 23799 18204 23811 18207
rect 24026 18204 24032 18216
rect 23799 18176 24032 18204
rect 23799 18173 23811 18176
rect 23753 18167 23811 18173
rect 24026 18164 24032 18176
rect 24084 18204 24090 18216
rect 24084 18176 24900 18204
rect 24084 18164 24090 18176
rect 19334 18136 19340 18148
rect 18524 18108 19340 18136
rect 19334 18096 19340 18108
rect 19392 18096 19398 18148
rect 22922 18096 22928 18148
rect 22980 18136 22986 18148
rect 24670 18136 24676 18148
rect 22980 18108 24676 18136
rect 22980 18096 22986 18108
rect 23860 18080 23888 18108
rect 24670 18096 24676 18108
rect 24728 18096 24734 18148
rect 14737 18071 14795 18077
rect 14737 18068 14749 18071
rect 13832 18040 14749 18068
rect 14737 18037 14749 18040
rect 14783 18037 14795 18071
rect 14737 18031 14795 18037
rect 15378 18028 15384 18080
rect 15436 18068 15442 18080
rect 16853 18071 16911 18077
rect 16853 18068 16865 18071
rect 15436 18040 16865 18068
rect 15436 18028 15442 18040
rect 16853 18037 16865 18040
rect 16899 18037 16911 18071
rect 16853 18031 16911 18037
rect 17957 18071 18015 18077
rect 17957 18037 17969 18071
rect 18003 18068 18015 18071
rect 18138 18068 18144 18080
rect 18003 18040 18144 18068
rect 18003 18037 18015 18040
rect 17957 18031 18015 18037
rect 18138 18028 18144 18040
rect 18196 18028 18202 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19521 18071 19579 18077
rect 19521 18068 19533 18071
rect 18656 18040 19533 18068
rect 18656 18028 18662 18040
rect 19521 18037 19533 18040
rect 19567 18037 19579 18071
rect 19521 18031 19579 18037
rect 23201 18071 23259 18077
rect 23201 18037 23213 18071
rect 23247 18068 23259 18071
rect 23290 18068 23296 18080
rect 23247 18040 23296 18068
rect 23247 18037 23259 18040
rect 23201 18031 23259 18037
rect 23290 18028 23296 18040
rect 23348 18028 23354 18080
rect 23842 18068 23848 18080
rect 23755 18040 23848 18068
rect 23842 18028 23848 18040
rect 23900 18028 23906 18080
rect 24026 18068 24032 18080
rect 23987 18040 24032 18068
rect 24026 18028 24032 18040
rect 24084 18028 24090 18080
rect 24872 18068 24900 18176
rect 26050 18164 26056 18216
rect 26108 18204 26114 18216
rect 26145 18207 26203 18213
rect 26145 18204 26157 18207
rect 26108 18176 26157 18204
rect 26108 18164 26114 18176
rect 26145 18173 26157 18176
rect 26191 18173 26203 18207
rect 26145 18167 26203 18173
rect 25314 18068 25320 18080
rect 24872 18040 25320 18068
rect 25314 18028 25320 18040
rect 25372 18028 25378 18080
rect 28994 18068 29000 18080
rect 28955 18040 29000 18068
rect 28994 18028 29000 18040
rect 29052 18028 29058 18080
rect 1104 17978 48852 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 48852 17978
rect 1104 17904 48852 17926
rect 7561 17867 7619 17873
rect 7561 17833 7573 17867
rect 7607 17864 7619 17867
rect 8294 17864 8300 17876
rect 7607 17836 8300 17864
rect 7607 17833 7619 17836
rect 7561 17827 7619 17833
rect 8294 17824 8300 17836
rect 8352 17824 8358 17876
rect 8389 17867 8447 17873
rect 8389 17833 8401 17867
rect 8435 17864 8447 17867
rect 8435 17836 9444 17864
rect 8435 17833 8447 17836
rect 8389 17827 8447 17833
rect 9306 17756 9312 17808
rect 9364 17756 9370 17808
rect 1397 17731 1455 17737
rect 1397 17697 1409 17731
rect 1443 17728 1455 17731
rect 1578 17728 1584 17740
rect 1443 17700 1584 17728
rect 1443 17697 1455 17700
rect 1397 17691 1455 17697
rect 1578 17688 1584 17700
rect 1636 17688 1642 17740
rect 2774 17688 2780 17740
rect 2832 17728 2838 17740
rect 2832 17700 2877 17728
rect 7208 17700 8340 17728
rect 2832 17688 2838 17700
rect 7208 17669 7236 17700
rect 7193 17663 7251 17669
rect 7193 17629 7205 17663
rect 7239 17629 7251 17663
rect 7193 17623 7251 17629
rect 7926 17620 7932 17672
rect 7984 17660 7990 17672
rect 8205 17663 8263 17669
rect 8205 17660 8217 17663
rect 7984 17632 8217 17660
rect 7984 17620 7990 17632
rect 8205 17629 8217 17632
rect 8251 17629 8263 17663
rect 8205 17623 8263 17629
rect 1581 17595 1639 17601
rect 1581 17561 1593 17595
rect 1627 17592 1639 17595
rect 2130 17592 2136 17604
rect 1627 17564 2136 17592
rect 1627 17561 1639 17564
rect 1581 17555 1639 17561
rect 2130 17552 2136 17564
rect 2188 17552 2194 17604
rect 7374 17592 7380 17604
rect 7335 17564 7380 17592
rect 7374 17552 7380 17564
rect 7432 17592 7438 17604
rect 8021 17595 8079 17601
rect 7432 17564 7972 17592
rect 7432 17552 7438 17564
rect 7944 17524 7972 17564
rect 8021 17561 8033 17595
rect 8067 17592 8079 17595
rect 8312 17592 8340 17700
rect 9324 17669 9352 17756
rect 9416 17669 9444 17836
rect 10870 17824 10876 17876
rect 10928 17864 10934 17876
rect 12069 17867 12127 17873
rect 12069 17864 12081 17867
rect 10928 17836 12081 17864
rect 10928 17824 10934 17836
rect 12069 17833 12081 17836
rect 12115 17833 12127 17867
rect 12069 17827 12127 17833
rect 13541 17867 13599 17873
rect 13541 17833 13553 17867
rect 13587 17864 13599 17867
rect 13998 17864 14004 17876
rect 13587 17836 14004 17864
rect 13587 17833 13599 17836
rect 13541 17827 13599 17833
rect 13998 17824 14004 17836
rect 14056 17824 14062 17876
rect 18049 17867 18107 17873
rect 18049 17833 18061 17867
rect 18095 17864 18107 17867
rect 20622 17864 20628 17876
rect 18095 17836 19012 17864
rect 20583 17836 20628 17864
rect 18095 17833 18107 17836
rect 18049 17827 18107 17833
rect 13170 17796 13176 17808
rect 12273 17768 13176 17796
rect 9217 17663 9275 17669
rect 9217 17629 9229 17663
rect 9263 17629 9275 17663
rect 9217 17623 9275 17629
rect 9309 17663 9367 17669
rect 9309 17629 9321 17663
rect 9355 17629 9367 17663
rect 9309 17623 9367 17629
rect 9401 17663 9459 17669
rect 9401 17629 9413 17663
rect 9447 17629 9459 17663
rect 9582 17660 9588 17672
rect 9543 17632 9588 17660
rect 9401 17623 9459 17629
rect 9232 17592 9260 17623
rect 9582 17620 9588 17632
rect 9640 17620 9646 17672
rect 10410 17620 10416 17672
rect 10468 17660 10474 17672
rect 10689 17663 10747 17669
rect 10689 17660 10701 17663
rect 10468 17632 10701 17660
rect 10468 17620 10474 17632
rect 10689 17629 10701 17632
rect 10735 17629 10747 17663
rect 10689 17623 10747 17629
rect 10956 17663 11014 17669
rect 10956 17629 10968 17663
rect 11002 17660 11014 17663
rect 11790 17660 11796 17672
rect 11002 17632 11796 17660
rect 11002 17629 11014 17632
rect 10956 17623 11014 17629
rect 9490 17592 9496 17604
rect 8067 17564 9168 17592
rect 9232 17564 9496 17592
rect 8067 17561 8079 17564
rect 8021 17555 8079 17561
rect 8754 17524 8760 17536
rect 7944 17496 8760 17524
rect 8754 17484 8760 17496
rect 8812 17484 8818 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 9140 17524 9168 17564
rect 9490 17552 9496 17564
rect 9548 17552 9554 17604
rect 10704 17592 10732 17623
rect 11790 17620 11796 17632
rect 11848 17620 11854 17672
rect 12273 17592 12301 17768
rect 13170 17756 13176 17768
rect 13228 17756 13234 17808
rect 13906 17756 13912 17808
rect 13964 17796 13970 17808
rect 16577 17799 16635 17805
rect 16577 17796 16589 17799
rect 13964 17768 16589 17796
rect 13964 17756 13970 17768
rect 16577 17765 16589 17768
rect 16623 17765 16635 17799
rect 17586 17796 17592 17808
rect 17547 17768 17592 17796
rect 16577 17759 16635 17765
rect 17586 17756 17592 17768
rect 17644 17756 17650 17808
rect 18506 17796 18512 17808
rect 17972 17768 18512 17796
rect 15289 17731 15347 17737
rect 15289 17728 15301 17731
rect 10704 17564 12301 17592
rect 12406 17700 15301 17728
rect 9214 17524 9220 17536
rect 9127 17496 9220 17524
rect 9214 17484 9220 17496
rect 9272 17524 9278 17536
rect 12406 17524 12434 17700
rect 12986 17620 12992 17672
rect 13044 17660 13050 17672
rect 13173 17663 13231 17669
rect 13173 17660 13185 17663
rect 13044 17632 13185 17660
rect 13044 17620 13050 17632
rect 13173 17629 13185 17632
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13262 17620 13268 17672
rect 13320 17660 13326 17672
rect 14200 17669 14228 17700
rect 15289 17697 15301 17700
rect 15335 17697 15347 17731
rect 15289 17691 15347 17697
rect 13357 17663 13415 17669
rect 13357 17660 13369 17663
rect 13320 17632 13369 17660
rect 13320 17620 13326 17632
rect 13357 17629 13369 17632
rect 13403 17629 13415 17663
rect 13357 17623 13415 17629
rect 14185 17663 14243 17669
rect 14185 17629 14197 17663
rect 14231 17629 14243 17663
rect 14185 17623 14243 17629
rect 15013 17663 15071 17669
rect 15013 17629 15025 17663
rect 15059 17660 15071 17663
rect 15746 17660 15752 17672
rect 15059 17632 15752 17660
rect 15059 17629 15071 17632
rect 15013 17623 15071 17629
rect 15746 17620 15752 17632
rect 15804 17620 15810 17672
rect 16393 17663 16451 17669
rect 16393 17629 16405 17663
rect 16439 17660 16451 17663
rect 17972 17660 18000 17768
rect 18506 17756 18512 17768
rect 18564 17756 18570 17808
rect 16439 17632 18000 17660
rect 18156 17700 18460 17728
rect 16439 17629 16451 17632
rect 16393 17623 16451 17629
rect 14366 17592 14372 17604
rect 14327 17564 14372 17592
rect 14366 17552 14372 17564
rect 14424 17552 14430 17604
rect 17405 17595 17463 17601
rect 17405 17561 17417 17595
rect 17451 17592 17463 17595
rect 17678 17592 17684 17604
rect 17451 17564 17684 17592
rect 17451 17561 17463 17564
rect 17405 17555 17463 17561
rect 17678 17552 17684 17564
rect 17736 17552 17742 17604
rect 9272 17496 12434 17524
rect 14553 17527 14611 17533
rect 9272 17484 9278 17496
rect 14553 17493 14565 17527
rect 14599 17524 14611 17527
rect 15470 17524 15476 17536
rect 14599 17496 15476 17524
rect 14599 17493 14611 17496
rect 14553 17487 14611 17493
rect 15470 17484 15476 17496
rect 15528 17484 15534 17536
rect 16758 17484 16764 17536
rect 16816 17524 16822 17536
rect 18156 17524 18184 17700
rect 18230 17620 18236 17672
rect 18288 17660 18294 17672
rect 18432 17669 18460 17700
rect 18325 17663 18383 17669
rect 18325 17660 18337 17663
rect 18288 17632 18337 17660
rect 18288 17620 18294 17632
rect 18325 17629 18337 17632
rect 18371 17629 18383 17663
rect 18325 17623 18383 17629
rect 18414 17663 18472 17669
rect 18414 17629 18426 17663
rect 18460 17629 18472 17663
rect 18414 17623 18472 17629
rect 18509 17663 18567 17669
rect 18509 17629 18521 17663
rect 18555 17629 18567 17663
rect 18509 17623 18567 17629
rect 18693 17663 18751 17669
rect 18693 17629 18705 17663
rect 18739 17629 18751 17663
rect 18984 17660 19012 17836
rect 20622 17824 20628 17836
rect 20680 17824 20686 17876
rect 22462 17864 22468 17876
rect 21652 17836 22468 17864
rect 19242 17728 19248 17740
rect 19203 17700 19248 17728
rect 19242 17688 19248 17700
rect 19300 17688 19306 17740
rect 19501 17663 19559 17669
rect 19501 17660 19513 17663
rect 18984 17632 19513 17660
rect 18693 17623 18751 17629
rect 19501 17629 19513 17632
rect 19547 17629 19559 17663
rect 20806 17660 20812 17672
rect 19501 17623 19559 17629
rect 19628 17632 20812 17660
rect 18524 17592 18552 17623
rect 18598 17592 18604 17604
rect 18524 17564 18604 17592
rect 18598 17552 18604 17564
rect 18656 17552 18662 17604
rect 18708 17592 18736 17623
rect 18782 17592 18788 17604
rect 18708 17564 18788 17592
rect 18782 17552 18788 17564
rect 18840 17552 18846 17604
rect 18414 17524 18420 17536
rect 16816 17496 18420 17524
rect 16816 17484 16822 17496
rect 18414 17484 18420 17496
rect 18472 17484 18478 17536
rect 18506 17484 18512 17536
rect 18564 17524 18570 17536
rect 19628 17524 19656 17632
rect 20806 17620 20812 17632
rect 20864 17620 20870 17672
rect 21652 17669 21680 17836
rect 22462 17824 22468 17836
rect 22520 17824 22526 17876
rect 23014 17824 23020 17876
rect 23072 17864 23078 17876
rect 24118 17864 24124 17876
rect 23072 17836 24124 17864
rect 23072 17824 23078 17836
rect 24118 17824 24124 17836
rect 24176 17824 24182 17876
rect 24765 17867 24823 17873
rect 24765 17833 24777 17867
rect 24811 17833 24823 17867
rect 24765 17827 24823 17833
rect 25685 17867 25743 17873
rect 25685 17833 25697 17867
rect 25731 17864 25743 17867
rect 26142 17864 26148 17876
rect 25731 17836 26148 17864
rect 25731 17833 25743 17836
rect 25685 17827 25743 17833
rect 21913 17799 21971 17805
rect 21913 17765 21925 17799
rect 21959 17796 21971 17799
rect 22557 17799 22615 17805
rect 22557 17796 22569 17799
rect 21959 17768 22569 17796
rect 21959 17765 21971 17768
rect 21913 17759 21971 17765
rect 22557 17765 22569 17768
rect 22603 17796 22615 17799
rect 22646 17796 22652 17808
rect 22603 17768 22652 17796
rect 22603 17765 22615 17768
rect 22557 17759 22615 17765
rect 22646 17756 22652 17768
rect 22704 17796 22710 17808
rect 23474 17796 23480 17808
rect 22704 17768 23480 17796
rect 22704 17756 22710 17768
rect 23474 17756 23480 17768
rect 23532 17756 23538 17808
rect 21775 17731 21833 17737
rect 21775 17697 21787 17731
rect 21821 17728 21833 17731
rect 22922 17728 22928 17740
rect 21821 17700 22928 17728
rect 21821 17697 21833 17700
rect 21775 17691 21833 17697
rect 22922 17688 22928 17700
rect 22980 17688 22986 17740
rect 23201 17731 23259 17737
rect 23382 17736 23388 17740
rect 23201 17697 23213 17731
rect 23247 17728 23259 17731
rect 23308 17728 23388 17736
rect 23247 17708 23388 17728
rect 23247 17700 23336 17708
rect 23247 17697 23259 17700
rect 23201 17691 23259 17697
rect 23382 17688 23388 17708
rect 23440 17688 23446 17740
rect 24780 17728 24808 17827
rect 26142 17824 26148 17836
rect 26200 17824 26206 17876
rect 26878 17824 26884 17876
rect 26936 17864 26942 17876
rect 29917 17867 29975 17873
rect 29917 17864 29929 17867
rect 26936 17836 29929 17864
rect 26936 17824 26942 17836
rect 29917 17833 29929 17836
rect 29963 17833 29975 17867
rect 29917 17827 29975 17833
rect 24946 17756 24952 17808
rect 25004 17796 25010 17808
rect 26053 17799 26111 17805
rect 26053 17796 26065 17799
rect 25004 17768 26065 17796
rect 25004 17756 25010 17768
rect 26053 17765 26065 17768
rect 26099 17796 26111 17799
rect 27249 17799 27307 17805
rect 27249 17796 27261 17799
rect 26099 17768 27261 17796
rect 26099 17765 26111 17768
rect 26053 17759 26111 17765
rect 27249 17765 27261 17768
rect 27295 17796 27307 17799
rect 28074 17796 28080 17808
rect 27295 17768 28080 17796
rect 27295 17765 27307 17768
rect 27249 17759 27307 17765
rect 28074 17756 28080 17768
rect 28132 17796 28138 17808
rect 28537 17799 28595 17805
rect 28537 17796 28549 17799
rect 28132 17768 28549 17796
rect 28132 17756 28138 17768
rect 28537 17765 28549 17768
rect 28583 17765 28595 17799
rect 28537 17759 28595 17765
rect 27709 17731 27767 17737
rect 27709 17728 27721 17731
rect 24780 17700 27721 17728
rect 27709 17697 27721 17700
rect 27755 17697 27767 17731
rect 27709 17691 27767 17697
rect 27801 17731 27859 17737
rect 27801 17697 27813 17731
rect 27847 17697 27859 17731
rect 27801 17691 27859 17697
rect 21637 17663 21695 17669
rect 21637 17629 21649 17663
rect 21683 17629 21695 17663
rect 21637 17623 21695 17629
rect 22094 17620 22100 17672
rect 22152 17660 22158 17672
rect 22152 17632 22197 17660
rect 22152 17620 22158 17632
rect 22462 17620 22468 17672
rect 22520 17660 22526 17672
rect 23017 17663 23075 17669
rect 22520 17632 22968 17660
rect 22520 17620 22526 17632
rect 20622 17552 20628 17604
rect 20680 17592 20686 17604
rect 22646 17592 22652 17604
rect 20680 17564 22652 17592
rect 20680 17552 20686 17564
rect 22646 17552 22652 17564
rect 22704 17552 22710 17604
rect 22940 17592 22968 17632
rect 23017 17629 23029 17663
rect 23063 17660 23075 17663
rect 23290 17660 23296 17672
rect 23063 17632 23296 17660
rect 23063 17629 23075 17632
rect 23017 17623 23075 17629
rect 23290 17620 23296 17632
rect 23348 17660 23354 17672
rect 24489 17663 24547 17669
rect 24489 17660 24501 17663
rect 23348 17632 24501 17660
rect 23348 17620 23354 17632
rect 24489 17629 24501 17632
rect 24535 17629 24547 17663
rect 24489 17623 24547 17629
rect 24673 17663 24731 17669
rect 24673 17629 24685 17663
rect 24719 17629 24731 17663
rect 24673 17623 24731 17629
rect 24765 17663 24823 17669
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 25130 17660 25136 17672
rect 24811 17632 25136 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 24578 17592 24584 17604
rect 22940 17564 24584 17592
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 18564 17496 19656 17524
rect 18564 17484 18570 17496
rect 20070 17484 20076 17536
rect 20128 17524 20134 17536
rect 20346 17524 20352 17536
rect 20128 17496 20352 17524
rect 20128 17484 20134 17496
rect 20346 17484 20352 17496
rect 20404 17484 20410 17536
rect 22097 17527 22155 17533
rect 22097 17493 22109 17527
rect 22143 17524 22155 17527
rect 22278 17524 22284 17536
rect 22143 17496 22284 17524
rect 22143 17493 22155 17496
rect 22097 17487 22155 17493
rect 22278 17484 22284 17496
rect 22336 17484 22342 17536
rect 22462 17484 22468 17536
rect 22520 17524 22526 17536
rect 22922 17524 22928 17536
rect 22520 17496 22928 17524
rect 22520 17484 22526 17496
rect 22922 17484 22928 17496
rect 22980 17484 22986 17536
rect 23014 17484 23020 17536
rect 23072 17524 23078 17536
rect 24688 17524 24716 17623
rect 25130 17620 25136 17632
rect 25188 17620 25194 17672
rect 25866 17660 25872 17672
rect 25827 17632 25872 17660
rect 25866 17620 25872 17632
rect 25924 17620 25930 17672
rect 26145 17663 26203 17669
rect 26145 17629 26157 17663
rect 26191 17660 26203 17663
rect 27430 17660 27436 17672
rect 26191 17632 27436 17660
rect 26191 17629 26203 17632
rect 26145 17623 26203 17629
rect 25314 17552 25320 17604
rect 25372 17592 25378 17604
rect 26160 17592 26188 17623
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 27614 17660 27620 17672
rect 27575 17632 27620 17660
rect 27614 17620 27620 17632
rect 27672 17620 27678 17672
rect 25372 17564 26188 17592
rect 25372 17552 25378 17564
rect 24946 17524 24952 17536
rect 23072 17496 24716 17524
rect 24907 17496 24952 17524
rect 23072 17484 23078 17496
rect 24946 17484 24952 17496
rect 25004 17484 25010 17536
rect 27632 17524 27660 17620
rect 27724 17592 27752 17691
rect 27816 17660 27844 17691
rect 27890 17688 27896 17740
rect 27948 17728 27954 17740
rect 28721 17731 28779 17737
rect 28721 17728 28733 17731
rect 27948 17700 28733 17728
rect 27948 17688 27954 17700
rect 28721 17697 28733 17700
rect 28767 17697 28779 17731
rect 28721 17691 28779 17697
rect 29178 17688 29184 17740
rect 29236 17728 29242 17740
rect 30006 17728 30012 17740
rect 29236 17700 30012 17728
rect 29236 17688 29242 17700
rect 30006 17688 30012 17700
rect 30064 17688 30070 17740
rect 28166 17660 28172 17672
rect 27816 17632 28172 17660
rect 28166 17620 28172 17632
rect 28224 17620 28230 17672
rect 28442 17660 28448 17672
rect 28403 17632 28448 17660
rect 28442 17620 28448 17632
rect 28500 17620 28506 17672
rect 29270 17620 29276 17672
rect 29328 17660 29334 17672
rect 29733 17663 29791 17669
rect 29733 17660 29745 17663
rect 29328 17632 29745 17660
rect 29328 17620 29334 17632
rect 29733 17629 29745 17632
rect 29779 17629 29791 17663
rect 29733 17623 29791 17629
rect 46290 17620 46296 17672
rect 46348 17660 46354 17672
rect 47673 17663 47731 17669
rect 47673 17660 47685 17663
rect 46348 17632 47685 17660
rect 46348 17620 46354 17632
rect 47673 17629 47685 17632
rect 47719 17629 47731 17663
rect 47673 17623 47731 17629
rect 28994 17592 29000 17604
rect 27724 17564 29000 17592
rect 28994 17552 29000 17564
rect 29052 17552 29058 17604
rect 28350 17524 28356 17536
rect 27632 17496 28356 17524
rect 28350 17484 28356 17496
rect 28408 17484 28414 17536
rect 28718 17524 28724 17536
rect 28679 17496 28724 17524
rect 28718 17484 28724 17496
rect 28776 17484 28782 17536
rect 29549 17527 29607 17533
rect 29549 17493 29561 17527
rect 29595 17524 29607 17527
rect 29822 17524 29828 17536
rect 29595 17496 29828 17524
rect 29595 17493 29607 17496
rect 29549 17487 29607 17493
rect 29822 17484 29828 17496
rect 29880 17484 29886 17536
rect 1104 17434 48852 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 48852 17434
rect 1104 17360 48852 17382
rect 7926 17280 7932 17332
rect 7984 17320 7990 17332
rect 9217 17323 9275 17329
rect 9217 17320 9229 17323
rect 7984 17292 9229 17320
rect 7984 17280 7990 17292
rect 9217 17289 9229 17292
rect 9263 17289 9275 17323
rect 9217 17283 9275 17289
rect 9306 17280 9312 17332
rect 9364 17320 9370 17332
rect 9364 17292 18552 17320
rect 9364 17280 9370 17292
rect 1581 17255 1639 17261
rect 1581 17221 1593 17255
rect 1627 17252 1639 17255
rect 2866 17252 2872 17264
rect 1627 17224 2872 17252
rect 1627 17221 1639 17224
rect 1581 17215 1639 17221
rect 2866 17212 2872 17224
rect 2924 17212 2930 17264
rect 7374 17252 7380 17264
rect 3712 17224 7380 17252
rect 3712 17193 3740 17224
rect 7374 17212 7380 17224
rect 7432 17212 7438 17264
rect 15562 17252 15568 17264
rect 15396 17224 15568 17252
rect 3697 17187 3755 17193
rect 3697 17153 3709 17187
rect 3743 17153 3755 17187
rect 7834 17184 7840 17196
rect 7795 17156 7840 17184
rect 3697 17147 3755 17153
rect 7834 17144 7840 17156
rect 7892 17144 7898 17196
rect 8104 17187 8162 17193
rect 8104 17153 8116 17187
rect 8150 17184 8162 17187
rect 8938 17184 8944 17196
rect 8150 17156 8944 17184
rect 8150 17153 8162 17156
rect 8104 17147 8162 17153
rect 8938 17144 8944 17156
rect 8996 17144 9002 17196
rect 13446 17193 13452 17196
rect 13440 17184 13452 17193
rect 13407 17156 13452 17184
rect 13440 17147 13452 17156
rect 13446 17144 13452 17147
rect 13504 17144 13510 17196
rect 15396 17193 15424 17224
rect 15562 17212 15568 17224
rect 15620 17212 15626 17264
rect 18414 17252 18420 17264
rect 18064 17224 18420 17252
rect 15289 17187 15347 17193
rect 15289 17153 15301 17187
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 1394 17116 1400 17128
rect 1355 17088 1400 17116
rect 1394 17076 1400 17088
rect 1452 17076 1458 17128
rect 2774 17076 2780 17128
rect 2832 17116 2838 17128
rect 3878 17116 3884 17128
rect 2832 17088 2877 17116
rect 3839 17088 3884 17116
rect 2832 17076 2838 17088
rect 3878 17076 3884 17088
rect 3936 17076 3942 17128
rect 4062 17076 4068 17128
rect 4120 17116 4126 17128
rect 4157 17119 4215 17125
rect 4157 17116 4169 17119
rect 4120 17088 4169 17116
rect 4120 17076 4126 17088
rect 4157 17085 4169 17088
rect 4203 17085 4215 17119
rect 13170 17116 13176 17128
rect 13131 17088 13176 17116
rect 4157 17079 4215 17085
rect 13170 17076 13176 17088
rect 13228 17076 13234 17128
rect 15010 17116 15016 17128
rect 14971 17088 15016 17116
rect 15010 17076 15016 17088
rect 15068 17076 15074 17128
rect 15304 17116 15332 17147
rect 15470 17144 15476 17196
rect 15528 17184 15534 17196
rect 15528 17156 15573 17184
rect 15528 17144 15534 17156
rect 15654 17144 15660 17196
rect 15712 17184 15718 17196
rect 16758 17184 16764 17196
rect 15712 17156 15757 17184
rect 16719 17156 16764 17184
rect 15712 17144 15718 17156
rect 16758 17144 16764 17156
rect 16816 17144 16822 17196
rect 16942 17184 16948 17196
rect 16903 17156 16948 17184
rect 16942 17144 16948 17156
rect 17000 17144 17006 17196
rect 17402 17184 17408 17196
rect 17363 17156 17408 17184
rect 17402 17144 17408 17156
rect 17460 17144 17466 17196
rect 17586 17184 17592 17196
rect 17547 17156 17592 17184
rect 17586 17144 17592 17156
rect 17644 17144 17650 17196
rect 18064 17193 18092 17224
rect 18414 17212 18420 17224
rect 18472 17212 18478 17264
rect 18524 17252 18552 17292
rect 18598 17280 18604 17332
rect 18656 17320 18662 17332
rect 19242 17320 19248 17332
rect 18656 17292 19248 17320
rect 18656 17280 18662 17292
rect 19242 17280 19248 17292
rect 19300 17320 19306 17332
rect 20257 17323 20315 17329
rect 20257 17320 20269 17323
rect 19300 17292 20269 17320
rect 19300 17280 19306 17292
rect 20257 17289 20269 17292
rect 20303 17289 20315 17323
rect 20257 17283 20315 17289
rect 22557 17323 22615 17329
rect 22557 17289 22569 17323
rect 22603 17320 22615 17323
rect 23477 17323 23535 17329
rect 23477 17320 23489 17323
rect 22603 17292 23489 17320
rect 22603 17289 22615 17292
rect 22557 17283 22615 17289
rect 23477 17289 23489 17292
rect 23523 17289 23535 17323
rect 23477 17283 23535 17289
rect 24854 17280 24860 17332
rect 24912 17320 24918 17332
rect 25133 17323 25191 17329
rect 25133 17320 25145 17323
rect 24912 17292 25145 17320
rect 24912 17280 24918 17292
rect 25133 17289 25145 17292
rect 25179 17289 25191 17323
rect 26326 17320 26332 17332
rect 26287 17292 26332 17320
rect 25133 17283 25191 17289
rect 26326 17280 26332 17292
rect 26384 17280 26390 17332
rect 30006 17320 30012 17332
rect 29967 17292 30012 17320
rect 30006 17280 30012 17292
rect 30064 17280 30070 17332
rect 23290 17252 23296 17264
rect 18524 17224 22876 17252
rect 18049 17187 18107 17193
rect 18049 17153 18061 17187
rect 18095 17153 18107 17187
rect 18049 17147 18107 17153
rect 18138 17144 18144 17196
rect 18196 17184 18202 17196
rect 18305 17187 18363 17193
rect 18305 17184 18317 17187
rect 18196 17156 18317 17184
rect 18196 17144 18202 17156
rect 18305 17153 18317 17156
rect 18351 17153 18363 17187
rect 18305 17147 18363 17153
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20165 17187 20223 17193
rect 20165 17184 20177 17187
rect 19668 17156 20177 17184
rect 19668 17144 19674 17156
rect 20165 17153 20177 17156
rect 20211 17153 20223 17187
rect 20165 17147 20223 17153
rect 21821 17187 21879 17193
rect 21821 17153 21833 17187
rect 21867 17184 21879 17187
rect 22462 17184 22468 17196
rect 21867 17156 22468 17184
rect 21867 17153 21879 17156
rect 21821 17147 21879 17153
rect 16574 17116 16580 17128
rect 15304 17088 16580 17116
rect 16574 17076 16580 17088
rect 16632 17076 16638 17128
rect 14550 17048 14556 17060
rect 14511 17020 14556 17048
rect 14550 17008 14556 17020
rect 14608 17008 14614 17060
rect 14826 17008 14832 17060
rect 14884 17048 14890 17060
rect 14884 17020 15056 17048
rect 14884 17008 14890 17020
rect 1762 16940 1768 16992
rect 1820 16980 1826 16992
rect 9306 16980 9312 16992
rect 1820 16952 9312 16980
rect 1820 16940 1826 16952
rect 9306 16940 9312 16952
rect 9364 16940 9370 16992
rect 15028 16980 15056 17020
rect 15102 17008 15108 17060
rect 15160 17048 15166 17060
rect 15654 17048 15660 17060
rect 15160 17020 15660 17048
rect 15160 17008 15166 17020
rect 15654 17008 15660 17020
rect 15712 17008 15718 17060
rect 19426 17048 19432 17060
rect 19339 17020 19432 17048
rect 19426 17008 19432 17020
rect 19484 17048 19490 17060
rect 21836 17048 21864 17147
rect 22462 17144 22468 17156
rect 22520 17144 22526 17196
rect 22097 17119 22155 17125
rect 22097 17085 22109 17119
rect 22143 17116 22155 17119
rect 22646 17116 22652 17128
rect 22143 17088 22652 17116
rect 22143 17085 22155 17088
rect 22097 17079 22155 17085
rect 22646 17076 22652 17088
rect 22704 17076 22710 17128
rect 22848 17116 22876 17224
rect 22940 17224 23296 17252
rect 22940 17193 22968 17224
rect 23290 17212 23296 17224
rect 23348 17212 23354 17264
rect 23382 17212 23388 17264
rect 23440 17252 23446 17264
rect 24673 17255 24731 17261
rect 24673 17252 24685 17255
rect 23440 17224 24685 17252
rect 23440 17212 23446 17224
rect 24673 17221 24685 17224
rect 24719 17221 24731 17255
rect 24673 17215 24731 17221
rect 27614 17212 27620 17264
rect 27672 17252 27678 17264
rect 28718 17252 28724 17264
rect 27672 17224 28724 17252
rect 27672 17212 27678 17224
rect 28718 17212 28724 17224
rect 28776 17212 28782 17264
rect 29089 17255 29147 17261
rect 29089 17221 29101 17255
rect 29135 17252 29147 17255
rect 29454 17252 29460 17264
rect 29135 17224 29460 17252
rect 29135 17221 29147 17224
rect 29089 17215 29147 17221
rect 29454 17212 29460 17224
rect 29512 17212 29518 17264
rect 31018 17212 31024 17264
rect 31076 17252 31082 17264
rect 46382 17252 46388 17264
rect 31076 17224 46388 17252
rect 31076 17212 31082 17224
rect 46382 17212 46388 17224
rect 46440 17212 46446 17264
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23017 17187 23075 17193
rect 23017 17153 23029 17187
rect 23063 17184 23075 17187
rect 23063 17156 23152 17184
rect 23063 17153 23075 17156
rect 23017 17147 23075 17153
rect 23124 17116 23152 17156
rect 23198 17144 23204 17196
rect 23256 17184 23262 17196
rect 23658 17184 23664 17196
rect 23256 17156 23301 17184
rect 23619 17156 23664 17184
rect 23256 17144 23262 17156
rect 23658 17144 23664 17156
rect 23716 17144 23722 17196
rect 23753 17187 23811 17193
rect 23753 17153 23765 17187
rect 23799 17184 23811 17187
rect 24026 17184 24032 17196
rect 23799 17156 24032 17184
rect 23799 17153 23811 17156
rect 23753 17147 23811 17153
rect 24026 17144 24032 17156
rect 24084 17144 24090 17196
rect 24949 17187 25007 17193
rect 24949 17184 24961 17187
rect 24136 17156 24961 17184
rect 22848 17088 23060 17116
rect 23124 17088 23336 17116
rect 19484 17020 21864 17048
rect 22005 17051 22063 17057
rect 19484 17008 19490 17020
rect 22005 17017 22017 17051
rect 22051 17048 22063 17051
rect 22462 17048 22468 17060
rect 22051 17020 22468 17048
rect 22051 17017 22063 17020
rect 22005 17011 22063 17017
rect 22462 17008 22468 17020
rect 22520 17008 22526 17060
rect 16853 16983 16911 16989
rect 16853 16980 16865 16983
rect 15028 16952 16865 16980
rect 16853 16949 16865 16952
rect 16899 16949 16911 16983
rect 16853 16943 16911 16949
rect 17497 16983 17555 16989
rect 17497 16949 17509 16983
rect 17543 16980 17555 16983
rect 18414 16980 18420 16992
rect 17543 16952 18420 16980
rect 17543 16949 17555 16952
rect 17497 16943 17555 16949
rect 18414 16940 18420 16952
rect 18472 16940 18478 16992
rect 18782 16940 18788 16992
rect 18840 16980 18846 16992
rect 20622 16980 20628 16992
rect 18840 16952 20628 16980
rect 18840 16940 18846 16952
rect 20622 16940 20628 16952
rect 20680 16940 20686 16992
rect 21913 16983 21971 16989
rect 21913 16949 21925 16983
rect 21959 16980 21971 16983
rect 22370 16980 22376 16992
rect 21959 16952 22376 16980
rect 21959 16949 21971 16952
rect 21913 16943 21971 16949
rect 22370 16940 22376 16952
rect 22428 16940 22434 16992
rect 23032 16980 23060 17088
rect 23308 17060 23336 17088
rect 23382 17076 23388 17128
rect 23440 17116 23446 17128
rect 23845 17119 23903 17125
rect 23845 17116 23857 17119
rect 23440 17088 23857 17116
rect 23440 17076 23446 17088
rect 23845 17085 23857 17088
rect 23891 17085 23903 17119
rect 23845 17079 23903 17085
rect 23937 17119 23995 17125
rect 23937 17085 23949 17119
rect 23983 17085 23995 17119
rect 23937 17079 23995 17085
rect 23290 17008 23296 17060
rect 23348 17008 23354 17060
rect 23658 17008 23664 17060
rect 23716 17048 23722 17060
rect 23952 17048 23980 17079
rect 23716 17020 23980 17048
rect 23716 17008 23722 17020
rect 24136 16980 24164 17156
rect 24949 17153 24961 17156
rect 24995 17153 25007 17187
rect 24949 17147 25007 17153
rect 26050 17144 26056 17196
rect 26108 17184 26114 17196
rect 26145 17187 26203 17193
rect 26145 17184 26157 17187
rect 26108 17156 26157 17184
rect 26108 17144 26114 17156
rect 26145 17153 26157 17156
rect 26191 17184 26203 17187
rect 28166 17184 28172 17196
rect 26191 17156 28172 17184
rect 26191 17153 26203 17156
rect 26145 17147 26203 17153
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 28902 17184 28908 17196
rect 28863 17156 28908 17184
rect 28902 17144 28908 17156
rect 28960 17144 28966 17196
rect 29178 17144 29184 17196
rect 29236 17184 29242 17196
rect 29236 17156 29281 17184
rect 29236 17144 29242 17156
rect 31662 17144 31668 17196
rect 31720 17184 31726 17196
rect 32125 17187 32183 17193
rect 32125 17184 32137 17187
rect 31720 17156 32137 17184
rect 31720 17144 31726 17156
rect 32125 17153 32137 17156
rect 32171 17153 32183 17187
rect 32125 17147 32183 17153
rect 32392 17187 32450 17193
rect 32392 17153 32404 17187
rect 32438 17184 32450 17187
rect 33502 17184 33508 17196
rect 32438 17156 33508 17184
rect 32438 17153 32450 17156
rect 32392 17147 32450 17153
rect 33502 17144 33508 17156
rect 33560 17144 33566 17196
rect 47210 17144 47216 17196
rect 47268 17184 47274 17196
rect 47581 17187 47639 17193
rect 47581 17184 47593 17187
rect 47268 17156 47593 17184
rect 47268 17144 47274 17156
rect 47581 17153 47593 17156
rect 47627 17153 47639 17187
rect 47581 17147 47639 17153
rect 24578 17076 24584 17128
rect 24636 17116 24642 17128
rect 24857 17119 24915 17125
rect 24636 17088 24808 17116
rect 24636 17076 24642 17088
rect 24210 17008 24216 17060
rect 24268 17048 24274 17060
rect 24780 17048 24808 17088
rect 24857 17085 24869 17119
rect 24903 17116 24915 17119
rect 25866 17116 25872 17128
rect 24903 17088 25872 17116
rect 24903 17085 24915 17088
rect 24857 17079 24915 17085
rect 25866 17076 25872 17088
rect 25924 17076 25930 17128
rect 27430 17116 27436 17128
rect 27391 17088 27436 17116
rect 27430 17076 27436 17088
rect 27488 17076 27494 17128
rect 27709 17119 27767 17125
rect 27709 17085 27721 17119
rect 27755 17116 27767 17119
rect 28442 17116 28448 17128
rect 27755 17088 28448 17116
rect 27755 17085 27767 17088
rect 27709 17079 27767 17085
rect 27724 17048 27752 17079
rect 28442 17076 28448 17088
rect 28500 17076 28506 17128
rect 30098 17116 30104 17128
rect 30059 17088 30104 17116
rect 30098 17076 30104 17088
rect 30156 17076 30162 17128
rect 30282 17116 30288 17128
rect 30243 17088 30288 17116
rect 30282 17076 30288 17088
rect 30340 17076 30346 17128
rect 24268 17020 24716 17048
rect 24780 17020 27752 17048
rect 28721 17051 28779 17057
rect 24268 17008 24274 17020
rect 24688 16989 24716 17020
rect 28721 17017 28733 17051
rect 28767 17048 28779 17051
rect 30006 17048 30012 17060
rect 28767 17020 30012 17048
rect 28767 17017 28779 17020
rect 28721 17011 28779 17017
rect 30006 17008 30012 17020
rect 30064 17008 30070 17060
rect 24305 16983 24363 16989
rect 24305 16980 24317 16983
rect 23032 16952 24317 16980
rect 24305 16949 24317 16952
rect 24351 16949 24363 16983
rect 24305 16943 24363 16949
rect 24673 16983 24731 16989
rect 24673 16949 24685 16983
rect 24719 16949 24731 16983
rect 24673 16943 24731 16949
rect 29178 16940 29184 16992
rect 29236 16980 29242 16992
rect 29641 16983 29699 16989
rect 29641 16980 29653 16983
rect 29236 16952 29653 16980
rect 29236 16940 29242 16952
rect 29641 16949 29653 16952
rect 29687 16949 29699 16983
rect 29641 16943 29699 16949
rect 29730 16940 29736 16992
rect 29788 16980 29794 16992
rect 32122 16980 32128 16992
rect 29788 16952 32128 16980
rect 29788 16940 29794 16952
rect 32122 16940 32128 16952
rect 32180 16940 32186 16992
rect 33042 16940 33048 16992
rect 33100 16980 33106 16992
rect 33505 16983 33563 16989
rect 33505 16980 33517 16983
rect 33100 16952 33517 16980
rect 33100 16940 33106 16952
rect 33505 16949 33517 16952
rect 33551 16949 33563 16983
rect 47026 16980 47032 16992
rect 46987 16952 47032 16980
rect 33505 16943 33563 16949
rect 47026 16940 47032 16952
rect 47084 16940 47090 16992
rect 47670 16980 47676 16992
rect 47631 16952 47676 16980
rect 47670 16940 47676 16952
rect 47728 16940 47734 16992
rect 1104 16890 48852 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 48852 16890
rect 1104 16816 48852 16838
rect 1394 16736 1400 16788
rect 1452 16776 1458 16788
rect 2685 16779 2743 16785
rect 2685 16776 2697 16779
rect 1452 16748 2697 16776
rect 1452 16736 1458 16748
rect 2685 16745 2697 16748
rect 2731 16745 2743 16779
rect 3878 16776 3884 16788
rect 3839 16748 3884 16776
rect 2685 16739 2743 16745
rect 3878 16736 3884 16748
rect 3936 16736 3942 16788
rect 7576 16748 16344 16776
rect 2041 16711 2099 16717
rect 2041 16677 2053 16711
rect 2087 16708 2099 16711
rect 7576 16708 7604 16748
rect 2087 16680 7604 16708
rect 2087 16677 2099 16680
rect 2041 16671 2099 16677
rect 13170 16668 13176 16720
rect 13228 16708 13234 16720
rect 13722 16708 13728 16720
rect 13228 16680 13728 16708
rect 13228 16668 13234 16680
rect 13722 16668 13728 16680
rect 13780 16708 13786 16720
rect 16316 16708 16344 16748
rect 16942 16736 16948 16788
rect 17000 16776 17006 16788
rect 17405 16779 17463 16785
rect 17405 16776 17417 16779
rect 17000 16748 17417 16776
rect 17000 16736 17006 16748
rect 17405 16745 17417 16748
rect 17451 16776 17463 16779
rect 17494 16776 17500 16788
rect 17451 16748 17500 16776
rect 17451 16745 17463 16748
rect 17405 16739 17463 16745
rect 17494 16736 17500 16748
rect 17552 16736 17558 16788
rect 17586 16736 17592 16788
rect 17644 16776 17650 16788
rect 17644 16748 18920 16776
rect 17644 16736 17650 16748
rect 18782 16708 18788 16720
rect 13780 16680 15424 16708
rect 16316 16680 18788 16708
rect 13780 16668 13786 16680
rect 15396 16652 15424 16680
rect 18782 16668 18788 16680
rect 18840 16668 18846 16720
rect 18892 16708 18920 16748
rect 19334 16736 19340 16788
rect 19392 16776 19398 16788
rect 19613 16779 19671 16785
rect 19613 16776 19625 16779
rect 19392 16748 19625 16776
rect 19392 16736 19398 16748
rect 19613 16745 19625 16748
rect 19659 16745 19671 16779
rect 19613 16739 19671 16745
rect 22646 16736 22652 16788
rect 22704 16776 22710 16788
rect 23661 16779 23719 16785
rect 22704 16748 23612 16776
rect 22704 16736 22710 16748
rect 20070 16708 20076 16720
rect 18892 16680 20076 16708
rect 20070 16668 20076 16680
rect 20128 16668 20134 16720
rect 22094 16668 22100 16720
rect 22152 16708 22158 16720
rect 23014 16708 23020 16720
rect 22152 16680 22416 16708
rect 22152 16668 22158 16680
rect 8018 16640 8024 16652
rect 3804 16612 8024 16640
rect 1854 16572 1860 16584
rect 1815 16544 1860 16572
rect 1854 16532 1860 16544
rect 1912 16532 1918 16584
rect 3804 16581 3832 16612
rect 8018 16600 8024 16612
rect 8076 16600 8082 16652
rect 10870 16600 10876 16652
rect 10928 16640 10934 16652
rect 10965 16643 11023 16649
rect 10965 16640 10977 16643
rect 10928 16612 10977 16640
rect 10928 16600 10934 16612
rect 10965 16609 10977 16612
rect 11011 16609 11023 16643
rect 11422 16640 11428 16652
rect 11383 16612 11428 16640
rect 10965 16603 11023 16609
rect 11422 16600 11428 16612
rect 11480 16600 11486 16652
rect 13906 16600 13912 16652
rect 13964 16640 13970 16652
rect 15378 16640 15384 16652
rect 13964 16612 14688 16640
rect 15339 16612 15384 16640
rect 13964 16600 13970 16612
rect 3789 16575 3847 16581
rect 3789 16541 3801 16575
rect 3835 16541 3847 16575
rect 14550 16572 14556 16584
rect 14511 16544 14556 16572
rect 3789 16535 3847 16541
rect 14550 16532 14556 16544
rect 14608 16532 14614 16584
rect 14660 16581 14688 16612
rect 15378 16600 15384 16612
rect 15436 16600 15442 16652
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 19610 16640 19616 16652
rect 19392 16612 19616 16640
rect 19392 16600 19398 16612
rect 19610 16600 19616 16612
rect 19668 16600 19674 16652
rect 22278 16600 22284 16652
rect 22336 16600 22342 16652
rect 14645 16575 14703 16581
rect 14645 16541 14657 16575
rect 14691 16541 14703 16575
rect 14645 16535 14703 16541
rect 14742 16575 14800 16581
rect 14742 16541 14754 16575
rect 14788 16574 14800 16575
rect 14921 16575 14979 16581
rect 14788 16546 14872 16574
rect 14788 16541 14800 16546
rect 14742 16535 14800 16541
rect 14844 16516 14872 16546
rect 14921 16541 14933 16575
rect 14967 16566 14979 16575
rect 15102 16566 15108 16584
rect 14967 16541 15108 16566
rect 14921 16538 15108 16541
rect 14921 16535 14979 16538
rect 15102 16532 15108 16538
rect 15160 16532 15166 16584
rect 17313 16575 17371 16581
rect 17313 16541 17325 16575
rect 17359 16572 17371 16575
rect 17586 16572 17592 16584
rect 17359 16544 17592 16572
rect 17359 16541 17371 16544
rect 17313 16535 17371 16541
rect 11149 16507 11207 16513
rect 11149 16473 11161 16507
rect 11195 16504 11207 16507
rect 11606 16504 11612 16516
rect 11195 16476 11612 16504
rect 11195 16473 11207 16476
rect 11149 16467 11207 16473
rect 11606 16464 11612 16476
rect 11664 16464 11670 16516
rect 14826 16464 14832 16516
rect 14884 16464 14890 16516
rect 15626 16507 15684 16513
rect 15626 16504 15638 16507
rect 14936 16476 15638 16504
rect 14 16396 20 16448
rect 72 16436 78 16448
rect 11422 16436 11428 16448
rect 72 16408 11428 16436
rect 72 16396 78 16408
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 14936 16436 14964 16476
rect 15626 16473 15638 16476
rect 15672 16473 15684 16507
rect 15626 16467 15684 16473
rect 14323 16408 14964 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 16574 16396 16580 16448
rect 16632 16436 16638 16448
rect 16761 16439 16819 16445
rect 16761 16436 16773 16439
rect 16632 16408 16773 16436
rect 16632 16396 16638 16408
rect 16761 16405 16773 16408
rect 16807 16436 16819 16439
rect 17328 16436 17356 16535
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 18509 16575 18567 16581
rect 18509 16541 18521 16575
rect 18555 16572 18567 16575
rect 20254 16572 20260 16584
rect 18555 16544 20260 16572
rect 18555 16541 18567 16544
rect 18509 16535 18567 16541
rect 20254 16532 20260 16544
rect 20312 16532 20318 16584
rect 20622 16572 20628 16584
rect 20583 16544 20628 16572
rect 20622 16532 20628 16544
rect 20680 16532 20686 16584
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 17678 16464 17684 16516
rect 17736 16504 17742 16516
rect 18690 16504 18696 16516
rect 17736 16476 18696 16504
rect 17736 16464 17742 16476
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 19245 16507 19303 16513
rect 19245 16473 19257 16507
rect 19291 16473 19303 16507
rect 19426 16504 19432 16516
rect 19387 16476 19432 16504
rect 19245 16467 19303 16473
rect 16807 16408 17356 16436
rect 19260 16436 19288 16467
rect 19426 16464 19432 16476
rect 19484 16464 19490 16516
rect 19518 16464 19524 16516
rect 19576 16464 19582 16516
rect 19536 16436 19564 16464
rect 22186 16436 22192 16448
rect 19260 16408 19564 16436
rect 22147 16408 22192 16436
rect 16807 16405 16819 16408
rect 16761 16399 16819 16405
rect 22186 16396 22192 16408
rect 22244 16396 22250 16448
rect 22296 16436 22324 16600
rect 22388 16572 22416 16680
rect 22664 16680 23020 16708
rect 22462 16600 22468 16652
rect 22520 16640 22526 16652
rect 22664 16649 22692 16680
rect 23014 16668 23020 16680
rect 23072 16668 23078 16720
rect 23584 16708 23612 16748
rect 23661 16745 23673 16779
rect 23707 16776 23719 16779
rect 23842 16776 23848 16788
rect 23707 16748 23848 16776
rect 23707 16745 23719 16748
rect 23661 16739 23719 16745
rect 23842 16736 23848 16748
rect 23900 16736 23906 16788
rect 25130 16736 25136 16788
rect 25188 16776 25194 16788
rect 25317 16779 25375 16785
rect 25317 16776 25329 16779
rect 25188 16748 25329 16776
rect 25188 16736 25194 16748
rect 25317 16745 25329 16748
rect 25363 16776 25375 16779
rect 25958 16776 25964 16788
rect 25363 16748 25964 16776
rect 25363 16745 25375 16748
rect 25317 16739 25375 16745
rect 25958 16736 25964 16748
rect 26016 16736 26022 16788
rect 28258 16776 28264 16788
rect 28219 16748 28264 16776
rect 28258 16736 28264 16748
rect 28316 16736 28322 16788
rect 31662 16776 31668 16788
rect 30944 16748 31668 16776
rect 24854 16708 24860 16720
rect 23584 16680 24860 16708
rect 24854 16668 24860 16680
rect 24912 16668 24918 16720
rect 28997 16711 29055 16717
rect 28997 16708 29009 16711
rect 27908 16680 29009 16708
rect 22649 16643 22707 16649
rect 22649 16640 22661 16643
rect 22520 16612 22661 16640
rect 22520 16600 22526 16612
rect 22649 16609 22661 16612
rect 22695 16609 22707 16643
rect 22649 16603 22707 16609
rect 22833 16643 22891 16649
rect 22833 16609 22845 16643
rect 22879 16640 22891 16643
rect 22922 16640 22928 16652
rect 22879 16612 22928 16640
rect 22879 16609 22891 16612
rect 22833 16603 22891 16609
rect 22922 16600 22928 16612
rect 22980 16600 22986 16652
rect 23474 16640 23480 16652
rect 23435 16612 23480 16640
rect 23474 16600 23480 16612
rect 23532 16600 23538 16652
rect 25869 16643 25927 16649
rect 25869 16609 25881 16643
rect 25915 16640 25927 16643
rect 26418 16640 26424 16652
rect 25915 16612 26424 16640
rect 25915 16609 25927 16612
rect 25869 16603 25927 16609
rect 26418 16600 26424 16612
rect 26476 16640 26482 16652
rect 27154 16640 27160 16652
rect 26476 16612 27160 16640
rect 26476 16600 26482 16612
rect 27154 16600 27160 16612
rect 27212 16600 27218 16652
rect 27908 16649 27936 16680
rect 28997 16677 29009 16680
rect 29043 16708 29055 16711
rect 29730 16708 29736 16720
rect 29043 16680 29736 16708
rect 29043 16677 29055 16680
rect 28997 16671 29055 16677
rect 29730 16668 29736 16680
rect 29788 16668 29794 16720
rect 30377 16711 30435 16717
rect 30377 16677 30389 16711
rect 30423 16708 30435 16711
rect 30742 16708 30748 16720
rect 30423 16680 30748 16708
rect 30423 16677 30435 16680
rect 30377 16671 30435 16677
rect 30742 16668 30748 16680
rect 30800 16668 30806 16720
rect 27893 16643 27951 16649
rect 27893 16609 27905 16643
rect 27939 16609 27951 16643
rect 29086 16640 29092 16652
rect 27893 16603 27951 16609
rect 28000 16612 29092 16640
rect 23385 16575 23443 16581
rect 23385 16572 23397 16575
rect 22388 16544 23397 16572
rect 23385 16541 23397 16544
rect 23431 16541 23443 16575
rect 23385 16535 23443 16541
rect 23661 16575 23719 16581
rect 23661 16541 23673 16575
rect 23707 16572 23719 16575
rect 25314 16572 25320 16584
rect 23707 16544 25320 16572
rect 23707 16541 23719 16544
rect 23661 16535 23719 16541
rect 25314 16532 25320 16544
rect 25372 16532 25378 16584
rect 26145 16575 26203 16581
rect 26145 16541 26157 16575
rect 26191 16541 26203 16575
rect 26145 16535 26203 16541
rect 22554 16504 22560 16516
rect 22467 16476 22560 16504
rect 22554 16464 22560 16476
rect 22612 16504 22618 16516
rect 23290 16504 23296 16516
rect 22612 16476 23296 16504
rect 22612 16464 22618 16476
rect 23290 16464 23296 16476
rect 23348 16464 23354 16516
rect 23474 16464 23480 16516
rect 23532 16504 23538 16516
rect 24486 16504 24492 16516
rect 23532 16476 24492 16504
rect 23532 16464 23538 16476
rect 24486 16464 24492 16476
rect 24544 16504 24550 16516
rect 25041 16507 25099 16513
rect 25041 16504 25053 16507
rect 24544 16476 25053 16504
rect 24544 16464 24550 16476
rect 25041 16473 25053 16476
rect 25087 16504 25099 16507
rect 26050 16504 26056 16516
rect 25087 16476 26056 16504
rect 25087 16473 25099 16476
rect 25041 16467 25099 16473
rect 26050 16464 26056 16476
rect 26108 16504 26114 16516
rect 26160 16504 26188 16535
rect 26970 16532 26976 16584
rect 27028 16572 27034 16584
rect 27246 16572 27252 16584
rect 27028 16544 27252 16572
rect 27028 16532 27034 16544
rect 27246 16532 27252 16544
rect 27304 16532 27310 16584
rect 27525 16575 27583 16581
rect 27525 16541 27537 16575
rect 27571 16572 27583 16575
rect 27614 16572 27620 16584
rect 27571 16544 27620 16572
rect 27571 16541 27583 16544
rect 27525 16535 27583 16541
rect 27614 16532 27620 16544
rect 27672 16532 27678 16584
rect 27709 16575 27767 16581
rect 27709 16541 27721 16575
rect 27755 16541 27767 16575
rect 27709 16535 27767 16541
rect 27801 16575 27859 16581
rect 27801 16541 27813 16575
rect 27847 16572 27859 16575
rect 28000 16572 28028 16612
rect 29086 16600 29092 16612
rect 29144 16600 29150 16652
rect 30944 16649 30972 16748
rect 31662 16736 31668 16748
rect 31720 16736 31726 16788
rect 33502 16776 33508 16788
rect 33463 16748 33508 16776
rect 33502 16736 33508 16748
rect 33560 16736 33566 16788
rect 32122 16668 32128 16720
rect 32180 16708 32186 16720
rect 32180 16680 33180 16708
rect 32180 16668 32186 16680
rect 30929 16643 30987 16649
rect 29656 16612 30144 16640
rect 27847 16544 28028 16572
rect 28077 16575 28135 16581
rect 27847 16541 27859 16544
rect 27801 16535 27859 16541
rect 28077 16541 28089 16575
rect 28123 16572 28135 16575
rect 28350 16572 28356 16584
rect 28123 16544 28356 16572
rect 28123 16541 28135 16544
rect 28077 16535 28135 16541
rect 26108 16476 26188 16504
rect 26108 16464 26114 16476
rect 22646 16436 22652 16448
rect 22296 16408 22652 16436
rect 22646 16396 22652 16408
rect 22704 16396 22710 16448
rect 23014 16396 23020 16448
rect 23072 16436 23078 16448
rect 23845 16439 23903 16445
rect 23845 16436 23857 16439
rect 23072 16408 23857 16436
rect 23072 16396 23078 16408
rect 23845 16405 23857 16408
rect 23891 16405 23903 16439
rect 23845 16399 23903 16405
rect 24394 16396 24400 16448
rect 24452 16436 24458 16448
rect 25682 16436 25688 16448
rect 24452 16408 25688 16436
rect 24452 16396 24458 16408
rect 25682 16396 25688 16408
rect 25740 16396 25746 16448
rect 26418 16396 26424 16448
rect 26476 16436 26482 16448
rect 27724 16436 27752 16535
rect 28350 16532 28356 16544
rect 28408 16532 28414 16584
rect 28718 16464 28724 16516
rect 28776 16504 28782 16516
rect 28813 16507 28871 16513
rect 28813 16504 28825 16507
rect 28776 16476 28825 16504
rect 28776 16464 28782 16476
rect 28813 16473 28825 16476
rect 28859 16473 28871 16507
rect 29656 16504 29684 16612
rect 29822 16572 29828 16584
rect 29783 16544 29828 16572
rect 29822 16532 29828 16544
rect 29880 16532 29886 16584
rect 30006 16572 30012 16584
rect 29967 16544 30012 16572
rect 30006 16532 30012 16544
rect 30064 16532 30070 16584
rect 30116 16572 30144 16612
rect 30929 16609 30941 16643
rect 30975 16609 30987 16643
rect 33042 16640 33048 16652
rect 33003 16612 33048 16640
rect 30929 16603 30987 16609
rect 33042 16600 33048 16612
rect 33100 16600 33106 16652
rect 33152 16649 33180 16680
rect 33137 16643 33195 16649
rect 33137 16609 33149 16643
rect 33183 16609 33195 16643
rect 46290 16640 46296 16652
rect 46251 16612 46296 16640
rect 33137 16603 33195 16609
rect 46290 16600 46296 16612
rect 46348 16600 46354 16652
rect 48130 16640 48136 16652
rect 48091 16612 48136 16640
rect 48130 16600 48136 16612
rect 48188 16600 48194 16652
rect 30193 16575 30251 16581
rect 30193 16572 30205 16575
rect 30116 16544 30205 16572
rect 30193 16541 30205 16544
rect 30239 16541 30251 16575
rect 30193 16535 30251 16541
rect 30668 16544 31340 16572
rect 29730 16504 29736 16516
rect 29656 16476 29736 16504
rect 28813 16467 28871 16473
rect 29730 16464 29736 16476
rect 29788 16464 29794 16516
rect 30098 16504 30104 16516
rect 30059 16476 30104 16504
rect 30098 16464 30104 16476
rect 30156 16504 30162 16516
rect 30668 16504 30696 16544
rect 30156 16476 30696 16504
rect 30156 16464 30162 16476
rect 30742 16464 30748 16516
rect 30800 16504 30806 16516
rect 31174 16507 31232 16513
rect 31174 16504 31186 16507
rect 30800 16476 31186 16504
rect 30800 16464 30806 16476
rect 31174 16473 31186 16476
rect 31220 16473 31232 16507
rect 31174 16467 31232 16473
rect 30926 16436 30932 16448
rect 26476 16408 30932 16436
rect 26476 16396 26482 16408
rect 30926 16396 30932 16408
rect 30984 16396 30990 16448
rect 31312 16436 31340 16544
rect 31570 16532 31576 16584
rect 31628 16572 31634 16584
rect 32769 16575 32827 16581
rect 32769 16572 32781 16575
rect 31628 16544 32781 16572
rect 31628 16532 31634 16544
rect 32769 16541 32781 16544
rect 32815 16541 32827 16575
rect 32950 16572 32956 16584
rect 32911 16544 32956 16572
rect 32769 16535 32827 16541
rect 32950 16532 32956 16544
rect 33008 16532 33014 16584
rect 33321 16575 33379 16581
rect 33321 16541 33333 16575
rect 33367 16541 33379 16575
rect 33321 16535 33379 16541
rect 31386 16464 31392 16516
rect 31444 16504 31450 16516
rect 33336 16504 33364 16535
rect 31444 16476 33364 16504
rect 46477 16507 46535 16513
rect 31444 16464 31450 16476
rect 46477 16473 46489 16507
rect 46523 16504 46535 16507
rect 47670 16504 47676 16516
rect 46523 16476 47676 16504
rect 46523 16473 46535 16476
rect 46477 16467 46535 16473
rect 47670 16464 47676 16476
rect 47728 16464 47734 16516
rect 32306 16436 32312 16448
rect 31312 16408 32312 16436
rect 32306 16396 32312 16408
rect 32364 16396 32370 16448
rect 1104 16346 48852 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 48852 16346
rect 1104 16272 48852 16294
rect 11606 16232 11612 16244
rect 11567 16204 11612 16232
rect 11606 16192 11612 16204
rect 11664 16192 11670 16244
rect 17494 16232 17500 16244
rect 17455 16204 17500 16232
rect 17494 16192 17500 16204
rect 17552 16192 17558 16244
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18693 16235 18751 16241
rect 18693 16232 18705 16235
rect 18472 16204 18705 16232
rect 18472 16192 18478 16204
rect 18693 16201 18705 16204
rect 18739 16201 18751 16235
rect 18693 16195 18751 16201
rect 21913 16235 21971 16241
rect 21913 16201 21925 16235
rect 21959 16232 21971 16235
rect 22094 16232 22100 16244
rect 21959 16204 22100 16232
rect 21959 16201 21971 16204
rect 21913 16195 21971 16201
rect 22094 16192 22100 16204
rect 22152 16192 22158 16244
rect 24394 16232 24400 16244
rect 23860 16204 24400 16232
rect 23860 16164 23888 16204
rect 24394 16192 24400 16204
rect 24452 16192 24458 16244
rect 28994 16232 29000 16244
rect 24596 16204 27016 16232
rect 28955 16204 29000 16232
rect 24026 16164 24032 16176
rect 12406 16136 23888 16164
rect 23939 16136 24032 16164
rect 11514 16096 11520 16108
rect 11475 16068 11520 16096
rect 11514 16056 11520 16068
rect 11572 16096 11578 16108
rect 12406 16096 12434 16136
rect 24026 16124 24032 16136
rect 24084 16164 24090 16176
rect 24596 16173 24624 16204
rect 24581 16167 24639 16173
rect 24581 16164 24593 16167
rect 24084 16136 24593 16164
rect 24084 16124 24090 16136
rect 24581 16133 24593 16136
rect 24627 16133 24639 16167
rect 24581 16127 24639 16133
rect 24670 16124 24676 16176
rect 24728 16164 24734 16176
rect 24765 16167 24823 16173
rect 24765 16164 24777 16167
rect 24728 16136 24777 16164
rect 24728 16124 24734 16136
rect 24765 16133 24777 16136
rect 24811 16133 24823 16167
rect 24765 16127 24823 16133
rect 24946 16124 24952 16176
rect 25004 16164 25010 16176
rect 25409 16167 25467 16173
rect 25409 16164 25421 16167
rect 25004 16136 25421 16164
rect 25004 16124 25010 16136
rect 25409 16133 25421 16136
rect 25455 16133 25467 16167
rect 25409 16127 25467 16133
rect 26988 16108 27016 16204
rect 28994 16192 29000 16204
rect 29052 16192 29058 16244
rect 30190 16232 30196 16244
rect 29380 16204 30196 16232
rect 27985 16167 28043 16173
rect 27985 16133 27997 16167
rect 28031 16164 28043 16167
rect 28442 16164 28448 16176
rect 28031 16136 28448 16164
rect 28031 16133 28043 16136
rect 27985 16127 28043 16133
rect 28442 16124 28448 16136
rect 28500 16124 28506 16176
rect 28629 16167 28687 16173
rect 28629 16133 28641 16167
rect 28675 16164 28687 16167
rect 29178 16164 29184 16176
rect 28675 16136 29184 16164
rect 28675 16133 28687 16136
rect 28629 16127 28687 16133
rect 29178 16124 29184 16136
rect 29236 16124 29242 16176
rect 13722 16096 13728 16108
rect 11572 16068 12434 16096
rect 13683 16068 13728 16096
rect 11572 16056 11578 16068
rect 13722 16056 13728 16068
rect 13780 16056 13786 16108
rect 13992 16099 14050 16105
rect 13992 16065 14004 16099
rect 14038 16096 14050 16099
rect 15010 16096 15016 16108
rect 14038 16068 15016 16096
rect 14038 16065 14050 16068
rect 13992 16059 14050 16065
rect 15010 16056 15016 16068
rect 15068 16056 15074 16108
rect 17310 16096 17316 16108
rect 17271 16068 17316 16096
rect 17310 16056 17316 16068
rect 17368 16056 17374 16108
rect 17402 16056 17408 16108
rect 17460 16096 17466 16108
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 17460 16068 17601 16096
rect 17460 16056 17466 16068
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 18509 16099 18567 16105
rect 18509 16096 18521 16099
rect 17589 16059 17647 16065
rect 18248 16068 18521 16096
rect 17328 16028 17356 16056
rect 17862 16028 17868 16040
rect 17328 16000 17868 16028
rect 17862 15988 17868 16000
rect 17920 16028 17926 16040
rect 18248 16028 18276 16068
rect 18509 16065 18521 16068
rect 18555 16065 18567 16099
rect 18782 16096 18788 16108
rect 18743 16068 18788 16096
rect 18509 16059 18567 16065
rect 18782 16056 18788 16068
rect 18840 16056 18846 16108
rect 19242 16096 19248 16108
rect 19203 16068 19248 16096
rect 19242 16056 19248 16068
rect 19300 16056 19306 16108
rect 19501 16099 19559 16105
rect 19501 16096 19513 16099
rect 19352 16068 19513 16096
rect 19352 16028 19380 16068
rect 19501 16065 19513 16068
rect 19547 16065 19559 16099
rect 19501 16059 19559 16065
rect 21821 16099 21879 16105
rect 21821 16065 21833 16099
rect 21867 16096 21879 16099
rect 22186 16096 22192 16108
rect 21867 16068 22192 16096
rect 21867 16065 21879 16068
rect 21821 16059 21879 16065
rect 22186 16056 22192 16068
rect 22244 16056 22250 16108
rect 22646 16096 22652 16108
rect 22607 16068 22652 16096
rect 22646 16056 22652 16068
rect 22704 16056 22710 16108
rect 22741 16099 22799 16105
rect 22741 16065 22753 16099
rect 22787 16096 22799 16099
rect 23014 16096 23020 16108
rect 22787 16068 23020 16096
rect 22787 16065 22799 16068
rect 22741 16059 22799 16065
rect 23014 16056 23020 16068
rect 23072 16056 23078 16108
rect 23658 16096 23664 16108
rect 23619 16068 23664 16096
rect 23658 16056 23664 16068
rect 23716 16056 23722 16108
rect 23845 16099 23903 16105
rect 23845 16065 23857 16099
rect 23891 16096 23903 16099
rect 23891 16068 24256 16096
rect 23891 16065 23903 16068
rect 23845 16059 23903 16065
rect 17920 16000 18276 16028
rect 18524 16000 19380 16028
rect 22833 16031 22891 16037
rect 17920 15988 17926 16000
rect 18524 15969 18552 16000
rect 22833 15997 22845 16031
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 18509 15963 18567 15969
rect 18509 15929 18521 15963
rect 18555 15929 18567 15963
rect 20622 15960 20628 15972
rect 20535 15932 20628 15960
rect 18509 15923 18567 15929
rect 20622 15920 20628 15932
rect 20680 15960 20686 15972
rect 22848 15960 22876 15991
rect 22922 15988 22928 16040
rect 22980 16028 22986 16040
rect 22980 16000 23025 16028
rect 22980 15988 22986 16000
rect 24118 15960 24124 15972
rect 20680 15932 22784 15960
rect 22848 15932 24124 15960
rect 20680 15920 20686 15932
rect 15102 15892 15108 15904
rect 15063 15864 15108 15892
rect 15102 15852 15108 15864
rect 15160 15852 15166 15904
rect 17126 15892 17132 15904
rect 17087 15864 17132 15892
rect 17126 15852 17132 15864
rect 17184 15852 17190 15904
rect 22278 15852 22284 15904
rect 22336 15892 22342 15904
rect 22465 15895 22523 15901
rect 22465 15892 22477 15895
rect 22336 15864 22477 15892
rect 22336 15852 22342 15864
rect 22465 15861 22477 15864
rect 22511 15861 22523 15895
rect 22756 15892 22784 15932
rect 24118 15920 24124 15932
rect 24176 15920 24182 15972
rect 24228 15960 24256 16068
rect 25038 16056 25044 16108
rect 25096 16096 25102 16108
rect 25685 16099 25743 16105
rect 25685 16096 25697 16099
rect 25096 16068 25697 16096
rect 25096 16056 25102 16068
rect 25685 16065 25697 16068
rect 25731 16065 25743 16099
rect 26970 16096 26976 16108
rect 26931 16068 26976 16096
rect 25685 16059 25743 16065
rect 26970 16056 26976 16068
rect 27028 16056 27034 16108
rect 27154 16096 27160 16108
rect 27115 16068 27160 16096
rect 27154 16056 27160 16068
rect 27212 16056 27218 16108
rect 27798 16096 27804 16108
rect 27759 16068 27804 16096
rect 27798 16056 27804 16068
rect 27856 16056 27862 16108
rect 28074 16096 28080 16108
rect 28035 16068 28080 16096
rect 28074 16056 28080 16068
rect 28132 16056 28138 16108
rect 28813 16099 28871 16105
rect 28813 16065 28825 16099
rect 28859 16096 28871 16099
rect 29380 16096 29408 16204
rect 30190 16192 30196 16204
rect 30248 16232 30254 16244
rect 30469 16235 30527 16241
rect 30469 16232 30481 16235
rect 30248 16204 30481 16232
rect 30248 16192 30254 16204
rect 30469 16201 30481 16204
rect 30515 16232 30527 16235
rect 30558 16232 30564 16244
rect 30515 16204 30564 16232
rect 30515 16201 30527 16204
rect 30469 16195 30527 16201
rect 30558 16192 30564 16204
rect 30616 16192 30622 16244
rect 30834 16164 30840 16176
rect 30795 16136 30840 16164
rect 30834 16124 30840 16136
rect 30892 16124 30898 16176
rect 30929 16167 30987 16173
rect 30929 16133 30941 16167
rect 30975 16164 30987 16167
rect 32125 16167 32183 16173
rect 32125 16164 32137 16167
rect 30975 16136 32137 16164
rect 30975 16133 30987 16136
rect 30929 16127 30987 16133
rect 32125 16133 32137 16136
rect 32171 16164 32183 16167
rect 33042 16164 33048 16176
rect 32171 16136 33048 16164
rect 32171 16133 32183 16136
rect 32125 16127 32183 16133
rect 33042 16124 33048 16136
rect 33100 16124 33106 16176
rect 28859 16068 29408 16096
rect 28859 16065 28871 16068
rect 28813 16059 28871 16065
rect 29454 16056 29460 16108
rect 29512 16096 29518 16108
rect 30852 16096 30880 16124
rect 31386 16096 31392 16108
rect 29512 16068 29557 16096
rect 30852 16068 31392 16096
rect 29512 16056 29518 16068
rect 31386 16056 31392 16068
rect 31444 16056 31450 16108
rect 32306 16096 32312 16108
rect 32267 16068 32312 16096
rect 32306 16056 32312 16068
rect 32364 16056 32370 16108
rect 32398 16056 32404 16108
rect 32456 16096 32462 16108
rect 32456 16068 32501 16096
rect 32456 16056 32462 16068
rect 47210 16056 47216 16108
rect 47268 16096 47274 16108
rect 47581 16099 47639 16105
rect 47581 16096 47593 16099
rect 47268 16068 47593 16096
rect 47268 16056 47274 16068
rect 47581 16065 47593 16068
rect 47627 16065 47639 16099
rect 47581 16059 47639 16065
rect 24854 15988 24860 16040
rect 24912 16028 24918 16040
rect 24949 16031 25007 16037
rect 24949 16028 24961 16031
rect 24912 16000 24961 16028
rect 24912 15988 24918 16000
rect 24949 15997 24961 16000
rect 24995 15997 25007 16031
rect 24949 15991 25007 15997
rect 25314 15988 25320 16040
rect 25372 16028 25378 16040
rect 25593 16031 25651 16037
rect 25593 16028 25605 16031
rect 25372 16000 25605 16028
rect 25372 15988 25378 16000
rect 25593 15997 25605 16000
rect 25639 16028 25651 16031
rect 29546 16028 29552 16040
rect 25639 16000 29552 16028
rect 25639 15997 25651 16000
rect 25593 15991 25651 15997
rect 29546 15988 29552 16000
rect 29604 15988 29610 16040
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 15997 29791 16031
rect 31018 16028 31024 16040
rect 30979 16000 31024 16028
rect 29733 15991 29791 15997
rect 25498 15960 25504 15972
rect 24228 15932 25504 15960
rect 24228 15892 24256 15932
rect 25498 15920 25504 15932
rect 25556 15920 25562 15972
rect 27801 15963 27859 15969
rect 27801 15929 27813 15963
rect 27847 15960 27859 15963
rect 27890 15960 27896 15972
rect 27847 15932 27896 15960
rect 27847 15929 27859 15932
rect 27801 15923 27859 15929
rect 27890 15920 27896 15932
rect 27948 15920 27954 15972
rect 29748 15960 29776 15991
rect 31018 15988 31024 16000
rect 31076 15988 31082 16040
rect 29196 15932 29776 15960
rect 30009 15963 30067 15969
rect 29196 15904 29224 15932
rect 30009 15929 30021 15963
rect 30055 15960 30067 15963
rect 30055 15932 31064 15960
rect 30055 15929 30067 15932
rect 30009 15923 30067 15929
rect 25590 15892 25596 15904
rect 22756 15864 24256 15892
rect 25551 15864 25596 15892
rect 22465 15855 22523 15861
rect 25590 15852 25596 15864
rect 25648 15852 25654 15904
rect 25869 15895 25927 15901
rect 25869 15861 25881 15895
rect 25915 15892 25927 15895
rect 26326 15892 26332 15904
rect 25915 15864 26332 15892
rect 25915 15861 25927 15864
rect 25869 15855 25927 15861
rect 26326 15852 26332 15864
rect 26384 15852 26390 15904
rect 27065 15895 27123 15901
rect 27065 15861 27077 15895
rect 27111 15892 27123 15895
rect 29178 15892 29184 15904
rect 27111 15864 29184 15892
rect 27111 15861 27123 15864
rect 27065 15855 27123 15861
rect 29178 15852 29184 15864
rect 29236 15852 29242 15904
rect 29825 15895 29883 15901
rect 29825 15861 29837 15895
rect 29871 15892 29883 15895
rect 30374 15892 30380 15904
rect 29871 15864 30380 15892
rect 29871 15861 29883 15864
rect 29825 15855 29883 15861
rect 30374 15852 30380 15864
rect 30432 15852 30438 15904
rect 31036 15892 31064 15932
rect 31570 15892 31576 15904
rect 31036 15864 31576 15892
rect 31570 15852 31576 15864
rect 31628 15852 31634 15904
rect 32122 15892 32128 15904
rect 32083 15864 32128 15892
rect 32122 15852 32128 15864
rect 32180 15852 32186 15904
rect 32306 15852 32312 15904
rect 32364 15892 32370 15904
rect 32585 15895 32643 15901
rect 32585 15892 32597 15895
rect 32364 15864 32597 15892
rect 32364 15852 32370 15864
rect 32585 15861 32597 15864
rect 32631 15861 32643 15895
rect 32585 15855 32643 15861
rect 46474 15852 46480 15904
rect 46532 15892 46538 15904
rect 47673 15895 47731 15901
rect 47673 15892 47685 15895
rect 46532 15864 47685 15892
rect 46532 15852 46538 15864
rect 47673 15861 47685 15864
rect 47719 15861 47731 15895
rect 47673 15855 47731 15861
rect 1104 15802 48852 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 48852 15802
rect 1104 15728 48852 15750
rect 17402 15648 17408 15700
rect 17460 15688 17466 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17460 15660 18153 15688
rect 17460 15648 17466 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 22462 15688 22468 15700
rect 22423 15660 22468 15688
rect 18141 15651 18199 15657
rect 22462 15648 22468 15660
rect 22520 15648 22526 15700
rect 22922 15688 22928 15700
rect 22883 15660 22928 15688
rect 22922 15648 22928 15660
rect 22980 15648 22986 15700
rect 24673 15691 24731 15697
rect 24673 15657 24685 15691
rect 24719 15688 24731 15691
rect 24762 15688 24768 15700
rect 24719 15660 24768 15688
rect 24719 15657 24731 15660
rect 24673 15651 24731 15657
rect 24762 15648 24768 15660
rect 24820 15648 24826 15700
rect 25501 15691 25559 15697
rect 25501 15657 25513 15691
rect 25547 15688 25559 15691
rect 25590 15688 25596 15700
rect 25547 15660 25596 15688
rect 25547 15657 25559 15660
rect 25501 15651 25559 15657
rect 25590 15648 25596 15660
rect 25648 15648 25654 15700
rect 26329 15691 26387 15697
rect 26329 15657 26341 15691
rect 26375 15688 26387 15691
rect 26970 15688 26976 15700
rect 26375 15660 26976 15688
rect 26375 15657 26387 15660
rect 26329 15651 26387 15657
rect 26970 15648 26976 15660
rect 27028 15648 27034 15700
rect 28629 15691 28687 15697
rect 28629 15657 28641 15691
rect 28675 15688 28687 15691
rect 28902 15688 28908 15700
rect 28675 15660 28908 15688
rect 28675 15657 28687 15660
rect 28629 15651 28687 15657
rect 28902 15648 28908 15660
rect 28960 15648 28966 15700
rect 30101 15691 30159 15697
rect 30101 15657 30113 15691
rect 30147 15657 30159 15691
rect 30101 15651 30159 15657
rect 14366 15620 14372 15632
rect 10612 15592 14372 15620
rect 10612 15561 10640 15592
rect 14366 15580 14372 15592
rect 14424 15620 14430 15632
rect 15102 15620 15108 15632
rect 14424 15592 15108 15620
rect 14424 15580 14430 15592
rect 15102 15580 15108 15592
rect 15160 15580 15166 15632
rect 17862 15580 17868 15632
rect 17920 15620 17926 15632
rect 19613 15623 19671 15629
rect 19613 15620 19625 15623
rect 17920 15592 19625 15620
rect 17920 15580 17926 15592
rect 19613 15589 19625 15592
rect 19659 15589 19671 15623
rect 25685 15623 25743 15629
rect 25685 15620 25697 15623
rect 19613 15583 19671 15589
rect 22103 15592 25697 15620
rect 10597 15555 10655 15561
rect 10597 15521 10609 15555
rect 10643 15521 10655 15555
rect 12342 15552 12348 15564
rect 12303 15524 12348 15552
rect 10597 15515 10655 15521
rect 12342 15512 12348 15524
rect 12400 15512 12406 15564
rect 19242 15512 19248 15564
rect 19300 15552 19306 15564
rect 21085 15555 21143 15561
rect 21085 15552 21097 15555
rect 19300 15524 21097 15552
rect 19300 15512 19306 15524
rect 21085 15521 21097 15524
rect 21131 15521 21143 15555
rect 21085 15515 21143 15521
rect 12894 15484 12900 15496
rect 12855 15456 12900 15484
rect 12894 15444 12900 15456
rect 12952 15444 12958 15496
rect 16761 15487 16819 15493
rect 16761 15453 16773 15487
rect 16807 15484 16819 15487
rect 19260 15484 19288 15512
rect 19426 15484 19432 15496
rect 16807 15456 19288 15484
rect 19387 15456 19432 15484
rect 16807 15453 16819 15456
rect 16761 15447 16819 15453
rect 19426 15444 19432 15456
rect 19484 15444 19490 15496
rect 22103 15484 22131 15592
rect 25685 15589 25697 15592
rect 25731 15589 25743 15623
rect 25685 15583 25743 15589
rect 28077 15623 28135 15629
rect 28077 15589 28089 15623
rect 28123 15620 28135 15623
rect 28166 15620 28172 15632
rect 28123 15592 28172 15620
rect 28123 15589 28135 15592
rect 28077 15583 28135 15589
rect 28166 15580 28172 15592
rect 28224 15620 28230 15632
rect 30006 15620 30012 15632
rect 28224 15592 30012 15620
rect 28224 15580 28230 15592
rect 30006 15580 30012 15592
rect 30064 15580 30070 15632
rect 25314 15552 25320 15564
rect 25275 15524 25320 15552
rect 25314 15512 25320 15524
rect 25372 15512 25378 15564
rect 26050 15512 26056 15564
rect 26108 15552 26114 15564
rect 30116 15552 30144 15651
rect 30282 15648 30288 15700
rect 30340 15688 30346 15700
rect 30837 15691 30895 15697
rect 30837 15688 30849 15691
rect 30340 15660 30849 15688
rect 30340 15648 30346 15660
rect 30837 15657 30849 15660
rect 30883 15657 30895 15691
rect 30837 15651 30895 15657
rect 30926 15580 30932 15632
rect 30984 15620 30990 15632
rect 31846 15620 31852 15632
rect 30984 15592 31852 15620
rect 30984 15580 30990 15592
rect 31846 15580 31852 15592
rect 31904 15620 31910 15632
rect 32950 15620 32956 15632
rect 31904 15592 32956 15620
rect 31904 15580 31910 15592
rect 26108 15524 27292 15552
rect 30116 15524 30558 15552
rect 26108 15512 26114 15524
rect 23106 15484 23112 15496
rect 21284 15456 22131 15484
rect 23067 15456 23112 15484
rect 10778 15416 10784 15428
rect 10739 15388 10784 15416
rect 10778 15376 10784 15388
rect 10836 15376 10842 15428
rect 17028 15419 17086 15425
rect 17028 15385 17040 15419
rect 17074 15416 17086 15419
rect 17126 15416 17132 15428
rect 17074 15388 17132 15416
rect 17074 15385 17086 15388
rect 17028 15379 17086 15385
rect 17126 15376 17132 15388
rect 17184 15376 17190 15428
rect 18782 15376 18788 15428
rect 18840 15416 18846 15428
rect 21284 15416 21312 15456
rect 23106 15444 23112 15456
rect 23164 15444 23170 15496
rect 23290 15484 23296 15496
rect 23251 15456 23296 15484
rect 23290 15444 23296 15456
rect 23348 15444 23354 15496
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15484 23443 15487
rect 24486 15484 24492 15496
rect 23431 15456 23520 15484
rect 24447 15456 24492 15484
rect 23431 15453 23443 15456
rect 23385 15447 23443 15453
rect 18840 15388 21312 15416
rect 21352 15419 21410 15425
rect 18840 15376 18846 15388
rect 21352 15385 21364 15419
rect 21398 15416 21410 15419
rect 22094 15416 22100 15428
rect 21398 15388 22100 15416
rect 21398 15385 21410 15388
rect 21352 15379 21410 15385
rect 22094 15376 22100 15388
rect 22152 15376 22158 15428
rect 12618 15308 12624 15360
rect 12676 15348 12682 15360
rect 13081 15351 13139 15357
rect 13081 15348 13093 15351
rect 12676 15320 13093 15348
rect 12676 15308 12682 15320
rect 13081 15317 13093 15320
rect 13127 15317 13139 15351
rect 13081 15311 13139 15317
rect 20990 15308 20996 15360
rect 21048 15348 21054 15360
rect 23492 15348 23520 15456
rect 24486 15444 24492 15456
rect 24544 15444 24550 15496
rect 24946 15444 24952 15496
rect 25004 15484 25010 15496
rect 25225 15487 25283 15493
rect 25225 15484 25237 15487
rect 25004 15456 25237 15484
rect 25004 15444 25010 15456
rect 25225 15453 25237 15456
rect 25271 15453 25283 15487
rect 25498 15484 25504 15496
rect 25459 15456 25504 15484
rect 25225 15447 25283 15453
rect 25498 15444 25504 15456
rect 25556 15444 25562 15496
rect 27065 15487 27123 15493
rect 27065 15453 27077 15487
rect 27111 15484 27123 15487
rect 27154 15484 27160 15496
rect 27111 15456 27160 15484
rect 27111 15453 27123 15456
rect 27065 15447 27123 15453
rect 27154 15444 27160 15456
rect 27212 15444 27218 15496
rect 27264 15484 27292 15524
rect 27264 15456 28396 15484
rect 24118 15376 24124 15428
rect 24176 15416 24182 15428
rect 26145 15419 26203 15425
rect 26145 15416 26157 15419
rect 24176 15388 26157 15416
rect 24176 15376 24182 15388
rect 26145 15385 26157 15388
rect 26191 15385 26203 15419
rect 26145 15379 26203 15385
rect 26326 15376 26332 15428
rect 26384 15425 26390 15428
rect 26384 15419 26403 15425
rect 26391 15385 26403 15419
rect 27890 15416 27896 15428
rect 27851 15388 27896 15416
rect 26384 15379 26403 15385
rect 26384 15376 26390 15379
rect 27890 15376 27896 15388
rect 27948 15376 27954 15428
rect 28368 15416 28396 15456
rect 28442 15444 28448 15496
rect 28500 15484 28506 15496
rect 28537 15487 28595 15493
rect 28537 15484 28549 15487
rect 28500 15456 28549 15484
rect 28500 15444 28506 15456
rect 28537 15453 28549 15456
rect 28583 15453 28595 15487
rect 28537 15447 28595 15453
rect 28718 15444 28724 15496
rect 28776 15484 28782 15496
rect 29825 15487 29883 15493
rect 28776 15456 28869 15484
rect 28776 15444 28782 15456
rect 29825 15453 29837 15487
rect 29871 15484 29883 15487
rect 30006 15484 30012 15496
rect 29871 15456 30012 15484
rect 29871 15453 29883 15456
rect 29825 15447 29883 15453
rect 30006 15444 30012 15456
rect 30064 15444 30070 15496
rect 30190 15484 30196 15496
rect 30151 15456 30196 15484
rect 30190 15444 30196 15456
rect 30248 15444 30254 15496
rect 30530 15484 30558 15524
rect 30742 15512 30748 15564
rect 30800 15552 30806 15564
rect 32140 15561 32168 15592
rect 32950 15580 32956 15592
rect 33008 15580 33014 15632
rect 47026 15620 47032 15632
rect 46308 15592 47032 15620
rect 46308 15561 46336 15592
rect 47026 15580 47032 15592
rect 47084 15580 47090 15632
rect 32033 15555 32091 15561
rect 32033 15552 32045 15555
rect 30800 15524 32045 15552
rect 30800 15512 30806 15524
rect 32033 15521 32045 15524
rect 32079 15521 32091 15555
rect 32033 15515 32091 15521
rect 32125 15555 32183 15561
rect 32125 15521 32137 15555
rect 32171 15521 32183 15555
rect 32125 15515 32183 15521
rect 46293 15555 46351 15561
rect 46293 15521 46305 15555
rect 46339 15521 46351 15555
rect 46474 15552 46480 15564
rect 46435 15524 46480 15552
rect 46293 15515 46351 15521
rect 46474 15512 46480 15524
rect 46532 15512 46538 15564
rect 48130 15552 48136 15564
rect 48091 15524 48136 15552
rect 48130 15512 48136 15524
rect 48188 15512 48194 15564
rect 30834 15484 30840 15496
rect 30530 15456 30840 15484
rect 30834 15444 30840 15456
rect 30892 15444 30898 15496
rect 30929 15487 30987 15493
rect 30929 15453 30941 15487
rect 30975 15453 30987 15487
rect 30929 15447 30987 15453
rect 28736 15416 28764 15444
rect 28368 15388 28764 15416
rect 29638 15376 29644 15428
rect 29696 15416 29702 15428
rect 30944 15416 30972 15447
rect 31754 15444 31760 15496
rect 31812 15484 31818 15496
rect 31812 15456 31857 15484
rect 31812 15444 31818 15456
rect 31938 15444 31944 15496
rect 31996 15484 32002 15496
rect 32309 15487 32367 15493
rect 31996 15456 32041 15484
rect 31996 15444 32002 15456
rect 32309 15453 32321 15487
rect 32355 15484 32367 15487
rect 32398 15484 32404 15496
rect 32355 15456 32404 15484
rect 32355 15453 32367 15456
rect 32309 15447 32367 15453
rect 32398 15444 32404 15456
rect 32456 15484 32462 15496
rect 33318 15484 33324 15496
rect 32456 15456 33324 15484
rect 32456 15444 32462 15456
rect 33318 15444 33324 15456
rect 33376 15484 33382 15496
rect 33962 15484 33968 15496
rect 33376 15456 33968 15484
rect 33376 15444 33382 15456
rect 33962 15444 33968 15456
rect 34020 15444 34026 15496
rect 29696 15388 30972 15416
rect 29696 15376 29702 15388
rect 26050 15348 26056 15360
rect 21048 15320 26056 15348
rect 21048 15308 21054 15320
rect 26050 15308 26056 15320
rect 26108 15308 26114 15360
rect 26510 15348 26516 15360
rect 26471 15320 26516 15348
rect 26510 15308 26516 15320
rect 26568 15308 26574 15360
rect 26878 15308 26884 15360
rect 26936 15348 26942 15360
rect 27157 15351 27215 15357
rect 27157 15348 27169 15351
rect 26936 15320 27169 15348
rect 26936 15308 26942 15320
rect 27157 15317 27169 15320
rect 27203 15317 27215 15351
rect 27157 15311 27215 15317
rect 29454 15308 29460 15360
rect 29512 15348 29518 15360
rect 30377 15351 30435 15357
rect 30377 15348 30389 15351
rect 29512 15320 30389 15348
rect 29512 15308 29518 15320
rect 30377 15317 30389 15320
rect 30423 15317 30435 15351
rect 30377 15311 30435 15317
rect 30466 15308 30472 15360
rect 30524 15348 30530 15360
rect 31205 15351 31263 15357
rect 31205 15348 31217 15351
rect 30524 15320 31217 15348
rect 30524 15308 30530 15320
rect 31205 15317 31217 15320
rect 31251 15317 31263 15351
rect 32490 15348 32496 15360
rect 32451 15320 32496 15348
rect 31205 15311 31263 15317
rect 32490 15308 32496 15320
rect 32548 15308 32554 15360
rect 1104 15258 48852 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 48852 15258
rect 1104 15184 48852 15206
rect 10778 15144 10784 15156
rect 10739 15116 10784 15144
rect 10778 15104 10784 15116
rect 10836 15104 10842 15156
rect 22094 15104 22100 15156
rect 22152 15144 22158 15156
rect 22152 15116 22197 15144
rect 22296 15116 24256 15144
rect 22152 15104 22158 15116
rect 22296 15076 22324 15116
rect 22066 15048 22324 15076
rect 10686 15008 10692 15020
rect 10647 14980 10692 15008
rect 10686 14968 10692 14980
rect 10744 14968 10750 15020
rect 19521 15011 19579 15017
rect 19521 14977 19533 15011
rect 19567 15008 19579 15011
rect 22066 15008 22094 15048
rect 23106 15036 23112 15088
rect 23164 15076 23170 15088
rect 23385 15079 23443 15085
rect 23385 15076 23397 15079
rect 23164 15048 23397 15076
rect 23164 15036 23170 15048
rect 23385 15045 23397 15048
rect 23431 15076 23443 15079
rect 24121 15079 24179 15085
rect 24121 15076 24133 15079
rect 23431 15048 24133 15076
rect 23431 15045 23443 15048
rect 23385 15039 23443 15045
rect 24121 15045 24133 15048
rect 24167 15045 24179 15079
rect 24121 15039 24179 15045
rect 22278 15008 22284 15020
rect 19567 14980 22094 15008
rect 22239 14980 22284 15008
rect 19567 14977 19579 14980
rect 19521 14971 19579 14977
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 22462 14968 22468 15020
rect 22520 15008 22526 15020
rect 22557 15011 22615 15017
rect 22557 15008 22569 15011
rect 22520 14980 22569 15008
rect 22520 14968 22526 14980
rect 22557 14977 22569 14980
rect 22603 14977 22615 15011
rect 24026 15008 24032 15020
rect 23987 14980 24032 15008
rect 22557 14971 22615 14977
rect 24026 14968 24032 14980
rect 24084 14968 24090 15020
rect 24228 15017 24256 15116
rect 25498 15104 25504 15156
rect 25556 15144 25562 15156
rect 25685 15147 25743 15153
rect 25685 15144 25697 15147
rect 25556 15116 25697 15144
rect 25556 15104 25562 15116
rect 25685 15113 25697 15116
rect 25731 15113 25743 15147
rect 25685 15107 25743 15113
rect 26237 15147 26295 15153
rect 26237 15113 26249 15147
rect 26283 15113 26295 15147
rect 26237 15107 26295 15113
rect 26252 15076 26280 15107
rect 27890 15104 27896 15156
rect 27948 15144 27954 15156
rect 28353 15147 28411 15153
rect 28353 15144 28365 15147
rect 27948 15116 28365 15144
rect 27948 15104 27954 15116
rect 28353 15113 28365 15116
rect 28399 15113 28411 15147
rect 29825 15147 29883 15153
rect 29825 15144 29837 15147
rect 28353 15107 28411 15113
rect 28460 15116 29837 15144
rect 27218 15079 27276 15085
rect 27218 15076 27230 15079
rect 26252 15048 27230 15076
rect 27218 15045 27230 15048
rect 27264 15045 27276 15079
rect 27218 15039 27276 15045
rect 27430 15036 27436 15088
rect 27488 15076 27494 15088
rect 28460 15076 28488 15116
rect 29825 15113 29837 15116
rect 29871 15113 29883 15147
rect 29825 15107 29883 15113
rect 30374 15104 30380 15156
rect 30432 15144 30438 15156
rect 30745 15147 30803 15153
rect 30745 15144 30757 15147
rect 30432 15116 30757 15144
rect 30432 15104 30438 15116
rect 30745 15113 30757 15116
rect 30791 15113 30803 15147
rect 30745 15107 30803 15113
rect 31573 15147 31631 15153
rect 31573 15113 31585 15147
rect 31619 15144 31631 15147
rect 31754 15144 31760 15156
rect 31619 15116 31760 15144
rect 31619 15113 31631 15116
rect 31573 15107 31631 15113
rect 31754 15104 31760 15116
rect 31812 15104 31818 15156
rect 33962 15144 33968 15156
rect 33923 15116 33968 15144
rect 33962 15104 33968 15116
rect 34020 15104 34026 15156
rect 46845 15147 46903 15153
rect 46845 15113 46857 15147
rect 46891 15144 46903 15147
rect 47854 15144 47860 15156
rect 46891 15116 47860 15144
rect 46891 15113 46903 15116
rect 46845 15107 46903 15113
rect 47854 15104 47860 15116
rect 47912 15104 47918 15156
rect 27488 15048 28488 15076
rect 27488 15036 27494 15048
rect 28994 15036 29000 15088
rect 29052 15076 29058 15088
rect 29365 15079 29423 15085
rect 29365 15076 29377 15079
rect 29052 15048 29377 15076
rect 29052 15036 29058 15048
rect 29365 15045 29377 15048
rect 29411 15045 29423 15079
rect 29365 15039 29423 15045
rect 29472 15048 30328 15076
rect 24213 15011 24271 15017
rect 24213 14977 24225 15011
rect 24259 15008 24271 15011
rect 24394 15008 24400 15020
rect 24259 14980 24400 15008
rect 24259 14977 24271 14980
rect 24213 14971 24271 14977
rect 24394 14968 24400 14980
rect 24452 15008 24458 15020
rect 24578 15008 24584 15020
rect 24452 14980 24584 15008
rect 24452 14968 24458 14980
rect 24578 14968 24584 14980
rect 24636 14968 24642 15020
rect 24765 15011 24823 15017
rect 24765 14977 24777 15011
rect 24811 15008 24823 15011
rect 24854 15008 24860 15020
rect 24811 14980 24860 15008
rect 24811 14977 24823 14980
rect 24765 14971 24823 14977
rect 24854 14968 24860 14980
rect 24912 14968 24918 15020
rect 25685 15011 25743 15017
rect 25685 14977 25697 15011
rect 25731 15008 25743 15011
rect 26142 15008 26148 15020
rect 25731 14980 26148 15008
rect 25731 14977 25743 14980
rect 25685 14971 25743 14977
rect 26142 14968 26148 14980
rect 26200 14968 26206 15020
rect 26421 15011 26479 15017
rect 26421 14977 26433 15011
rect 26467 15008 26479 15011
rect 26510 15008 26516 15020
rect 26467 14980 26516 15008
rect 26467 14977 26479 14980
rect 26421 14971 26479 14977
rect 26510 14968 26516 14980
rect 26568 14968 26574 15020
rect 27522 14968 27528 15020
rect 27580 15008 27586 15020
rect 29472 15008 29500 15048
rect 29638 15008 29644 15020
rect 27580 14980 29500 15008
rect 29599 14980 29644 15008
rect 27580 14968 27586 14980
rect 29638 14968 29644 14980
rect 29696 14968 29702 15020
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 19705 14943 19763 14949
rect 19705 14940 19717 14943
rect 19484 14912 19717 14940
rect 19484 14900 19490 14912
rect 19705 14909 19717 14912
rect 19751 14940 19763 14943
rect 20990 14940 20996 14952
rect 19751 14912 20996 14940
rect 19751 14909 19763 14912
rect 19705 14903 19763 14909
rect 20990 14900 20996 14912
rect 21048 14900 21054 14952
rect 26234 14900 26240 14952
rect 26292 14940 26298 14952
rect 26973 14943 27031 14949
rect 26973 14940 26985 14943
rect 26292 14912 26985 14940
rect 26292 14900 26298 14912
rect 26973 14909 26985 14912
rect 27019 14909 27031 14943
rect 29546 14940 29552 14952
rect 29507 14912 29552 14940
rect 26973 14903 27031 14909
rect 29546 14900 29552 14912
rect 29604 14900 29610 14952
rect 30300 14940 30328 15048
rect 32490 15036 32496 15088
rect 32548 15076 32554 15088
rect 32830 15079 32888 15085
rect 32830 15076 32842 15079
rect 32548 15048 32842 15076
rect 32548 15036 32554 15048
rect 32830 15045 32842 15048
rect 32876 15045 32888 15079
rect 32830 15039 32888 15045
rect 30466 15008 30472 15020
rect 30427 14980 30472 15008
rect 30466 14968 30472 14980
rect 30524 14968 30530 15020
rect 30558 14968 30564 15020
rect 30616 15008 30622 15020
rect 30616 14980 30661 15008
rect 30616 14968 30622 14980
rect 31018 14968 31024 15020
rect 31076 15008 31082 15020
rect 31205 15011 31263 15017
rect 31205 15008 31217 15011
rect 31076 14980 31217 15008
rect 31076 14968 31082 14980
rect 31205 14977 31217 14980
rect 31251 14977 31263 15011
rect 31205 14971 31263 14977
rect 31389 15011 31447 15017
rect 31389 14977 31401 15011
rect 31435 15008 31447 15011
rect 33226 15008 33232 15020
rect 31435 14980 33232 15008
rect 31435 14977 31447 14980
rect 31389 14971 31447 14977
rect 33226 14968 33232 14980
rect 33284 15008 33290 15020
rect 33870 15008 33876 15020
rect 33284 14980 33876 15008
rect 33284 14968 33290 14980
rect 33870 14968 33876 14980
rect 33928 14968 33934 15020
rect 46842 14968 46848 15020
rect 46900 15008 46906 15020
rect 47029 15011 47087 15017
rect 47029 15008 47041 15011
rect 46900 14980 47041 15008
rect 46900 14968 46906 14980
rect 47029 14977 47041 14980
rect 47075 14977 47087 15011
rect 47029 14971 47087 14977
rect 30300 14912 31754 14940
rect 15746 14832 15752 14884
rect 15804 14872 15810 14884
rect 18230 14872 18236 14884
rect 15804 14844 18236 14872
rect 15804 14832 15810 14844
rect 18230 14832 18236 14844
rect 18288 14872 18294 14884
rect 22465 14875 22523 14881
rect 18288 14844 22094 14872
rect 18288 14832 18294 14844
rect 22066 14804 22094 14844
rect 22465 14841 22477 14875
rect 22511 14872 22523 14875
rect 24762 14872 24768 14884
rect 22511 14844 24768 14872
rect 22511 14841 22523 14844
rect 22465 14835 22523 14841
rect 24762 14832 24768 14844
rect 24820 14832 24826 14884
rect 26878 14872 26884 14884
rect 24872 14844 26884 14872
rect 23382 14804 23388 14816
rect 22066 14776 23388 14804
rect 23382 14764 23388 14776
rect 23440 14764 23446 14816
rect 23474 14764 23480 14816
rect 23532 14804 23538 14816
rect 23658 14804 23664 14816
rect 23532 14776 23664 14804
rect 23532 14764 23538 14776
rect 23658 14764 23664 14776
rect 23716 14764 23722 14816
rect 23842 14764 23848 14816
rect 23900 14804 23906 14816
rect 24872 14804 24900 14844
rect 26878 14832 26884 14844
rect 26936 14832 26942 14884
rect 30282 14872 30288 14884
rect 29656 14844 30288 14872
rect 23900 14776 24900 14804
rect 24949 14807 25007 14813
rect 23900 14764 23906 14776
rect 24949 14773 24961 14807
rect 24995 14804 25007 14807
rect 25038 14804 25044 14816
rect 24995 14776 25044 14804
rect 24995 14773 25007 14776
rect 24949 14767 25007 14773
rect 25038 14764 25044 14776
rect 25096 14764 25102 14816
rect 26896 14804 26924 14832
rect 29362 14804 29368 14816
rect 26896 14776 29368 14804
rect 29362 14764 29368 14776
rect 29420 14764 29426 14816
rect 29454 14764 29460 14816
rect 29512 14804 29518 14816
rect 29656 14813 29684 14844
rect 30282 14832 30288 14844
rect 30340 14832 30346 14884
rect 31726 14872 31754 14912
rect 32398 14900 32404 14952
rect 32456 14940 32462 14952
rect 32585 14943 32643 14949
rect 32585 14940 32597 14943
rect 32456 14912 32597 14940
rect 32456 14900 32462 14912
rect 32585 14909 32597 14912
rect 32631 14909 32643 14943
rect 32585 14903 32643 14909
rect 32490 14872 32496 14884
rect 31726 14844 32496 14872
rect 32490 14832 32496 14844
rect 32548 14832 32554 14884
rect 29641 14807 29699 14813
rect 29641 14804 29653 14807
rect 29512 14776 29653 14804
rect 29512 14764 29518 14776
rect 29641 14773 29653 14776
rect 29687 14773 29699 14807
rect 47762 14804 47768 14816
rect 47723 14776 47768 14804
rect 29641 14767 29699 14773
rect 47762 14764 47768 14776
rect 47820 14764 47826 14816
rect 1104 14714 48852 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 48852 14714
rect 1104 14640 48852 14662
rect 19334 14560 19340 14612
rect 19392 14600 19398 14612
rect 19429 14603 19487 14609
rect 19429 14600 19441 14603
rect 19392 14572 19441 14600
rect 19392 14560 19398 14572
rect 19429 14569 19441 14572
rect 19475 14569 19487 14603
rect 19429 14563 19487 14569
rect 20254 14560 20260 14612
rect 20312 14600 20318 14612
rect 20312 14572 23060 14600
rect 20312 14560 20318 14572
rect 21269 14535 21327 14541
rect 21269 14501 21281 14535
rect 21315 14532 21327 14535
rect 21450 14532 21456 14544
rect 21315 14504 21456 14532
rect 21315 14501 21327 14504
rect 21269 14495 21327 14501
rect 21450 14492 21456 14504
rect 21508 14532 21514 14544
rect 21726 14532 21732 14544
rect 21508 14504 21732 14532
rect 21508 14492 21514 14504
rect 21726 14492 21732 14504
rect 21784 14492 21790 14544
rect 1762 14356 1768 14408
rect 1820 14396 1826 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1820 14368 2053 14396
rect 1820 14356 1826 14368
rect 2041 14365 2053 14368
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 18690 14356 18696 14408
rect 18748 14396 18754 14408
rect 19337 14399 19395 14405
rect 19337 14396 19349 14399
rect 18748 14368 19349 14396
rect 18748 14356 18754 14368
rect 19337 14365 19349 14368
rect 19383 14365 19395 14399
rect 19337 14359 19395 14365
rect 20806 14356 20812 14408
rect 20864 14396 20870 14408
rect 21085 14399 21143 14405
rect 21085 14396 21097 14399
rect 20864 14368 21097 14396
rect 20864 14356 20870 14368
rect 21085 14365 21097 14368
rect 21131 14365 21143 14399
rect 22830 14396 22836 14408
rect 22791 14368 22836 14396
rect 21085 14359 21143 14365
rect 22830 14356 22836 14368
rect 22888 14356 22894 14408
rect 23032 14405 23060 14572
rect 23474 14560 23480 14612
rect 23532 14600 23538 14612
rect 24486 14600 24492 14612
rect 23532 14572 24492 14600
rect 23532 14560 23538 14572
rect 24486 14560 24492 14572
rect 24544 14560 24550 14612
rect 25225 14603 25283 14609
rect 25225 14569 25237 14603
rect 25271 14600 25283 14603
rect 26418 14600 26424 14612
rect 25271 14572 26424 14600
rect 25271 14569 25283 14572
rect 25225 14563 25283 14569
rect 26418 14560 26424 14572
rect 26476 14560 26482 14612
rect 29546 14560 29552 14612
rect 29604 14600 29610 14612
rect 30193 14603 30251 14609
rect 30193 14600 30205 14603
rect 29604 14572 30205 14600
rect 29604 14560 29610 14572
rect 30193 14569 30205 14572
rect 30239 14600 30251 14603
rect 30834 14600 30840 14612
rect 30239 14572 30840 14600
rect 30239 14569 30251 14572
rect 30193 14563 30251 14569
rect 30834 14560 30840 14572
rect 30892 14560 30898 14612
rect 31205 14603 31263 14609
rect 31205 14569 31217 14603
rect 31251 14600 31263 14603
rect 31938 14600 31944 14612
rect 31251 14572 31944 14600
rect 31251 14569 31263 14572
rect 31205 14563 31263 14569
rect 31938 14560 31944 14572
rect 31996 14560 32002 14612
rect 32490 14560 32496 14612
rect 32548 14600 32554 14612
rect 48038 14600 48044 14612
rect 32548 14572 48044 14600
rect 32548 14560 32554 14572
rect 48038 14560 48044 14572
rect 48096 14560 48102 14612
rect 24762 14492 24768 14544
rect 24820 14532 24826 14544
rect 28905 14535 28963 14541
rect 28905 14532 28917 14535
rect 24820 14504 28917 14532
rect 24820 14492 24826 14504
rect 28905 14501 28917 14504
rect 28951 14501 28963 14535
rect 28905 14495 28963 14501
rect 29362 14492 29368 14544
rect 29420 14532 29426 14544
rect 31018 14532 31024 14544
rect 29420 14504 31024 14532
rect 29420 14492 29426 14504
rect 31018 14492 31024 14504
rect 31076 14492 31082 14544
rect 32861 14535 32919 14541
rect 32861 14532 32873 14535
rect 31726 14504 32873 14532
rect 25038 14424 25044 14476
rect 25096 14464 25102 14476
rect 30745 14467 30803 14473
rect 30745 14464 30757 14467
rect 25096 14436 28764 14464
rect 25096 14424 25102 14436
rect 23017 14399 23075 14405
rect 23017 14365 23029 14399
rect 23063 14396 23075 14399
rect 26605 14399 26663 14405
rect 26605 14396 26617 14399
rect 23063 14368 26617 14396
rect 23063 14365 23075 14368
rect 23017 14359 23075 14365
rect 26605 14365 26617 14368
rect 26651 14365 26663 14399
rect 26605 14359 26663 14365
rect 26789 14399 26847 14405
rect 26789 14365 26801 14399
rect 26835 14396 26847 14399
rect 27617 14399 27675 14405
rect 27617 14396 27629 14399
rect 26835 14368 27629 14396
rect 26835 14365 26847 14368
rect 26789 14359 26847 14365
rect 27617 14365 27629 14368
rect 27663 14396 27675 14399
rect 27982 14396 27988 14408
rect 27663 14368 27988 14396
rect 27663 14365 27675 14368
rect 27617 14359 27675 14365
rect 27982 14356 27988 14368
rect 28040 14356 28046 14408
rect 28736 14405 28764 14436
rect 29840 14436 30757 14464
rect 28721 14399 28779 14405
rect 28721 14365 28733 14399
rect 28767 14396 28779 14399
rect 29270 14396 29276 14408
rect 28767 14368 29276 14396
rect 28767 14365 28779 14368
rect 28721 14359 28779 14365
rect 29270 14356 29276 14368
rect 29328 14356 29334 14408
rect 29840 14405 29868 14436
rect 30745 14433 30757 14436
rect 30791 14464 30803 14467
rect 31726 14464 31754 14504
rect 32861 14501 32873 14504
rect 32907 14501 32919 14535
rect 32861 14495 32919 14501
rect 30791 14436 31754 14464
rect 31941 14467 31999 14473
rect 30791 14433 30803 14436
rect 30745 14427 30803 14433
rect 31941 14433 31953 14467
rect 31987 14464 31999 14467
rect 32122 14464 32128 14476
rect 31987 14436 32128 14464
rect 31987 14433 31999 14436
rect 31941 14427 31999 14433
rect 32122 14424 32128 14436
rect 32180 14424 32186 14476
rect 33318 14464 33324 14476
rect 33279 14436 33324 14464
rect 33318 14424 33324 14436
rect 33376 14424 33382 14476
rect 33413 14467 33471 14473
rect 33413 14433 33425 14467
rect 33459 14433 33471 14467
rect 33413 14427 33471 14433
rect 46293 14467 46351 14473
rect 46293 14433 46305 14467
rect 46339 14464 46351 14467
rect 47762 14464 47768 14476
rect 46339 14436 47768 14464
rect 46339 14433 46351 14436
rect 46293 14427 46351 14433
rect 29825 14399 29883 14405
rect 29825 14365 29837 14399
rect 29871 14365 29883 14399
rect 30558 14396 30564 14408
rect 29825 14359 29883 14365
rect 29932 14368 30564 14396
rect 20257 14331 20315 14337
rect 20257 14297 20269 14331
rect 20303 14328 20315 14331
rect 24670 14328 24676 14340
rect 20303 14300 24676 14328
rect 20303 14297 20315 14300
rect 20257 14291 20315 14297
rect 24670 14288 24676 14300
rect 24728 14288 24734 14340
rect 24854 14288 24860 14340
rect 24912 14328 24918 14340
rect 25133 14331 25191 14337
rect 25133 14328 25145 14331
rect 24912 14300 25145 14328
rect 24912 14288 24918 14300
rect 25133 14297 25145 14300
rect 25179 14297 25191 14331
rect 27798 14328 27804 14340
rect 27759 14300 27804 14328
rect 25133 14291 25191 14297
rect 27798 14288 27804 14300
rect 27856 14288 27862 14340
rect 20533 14263 20591 14269
rect 20533 14229 20545 14263
rect 20579 14260 20591 14263
rect 21174 14260 21180 14272
rect 20579 14232 21180 14260
rect 20579 14229 20591 14232
rect 20533 14223 20591 14229
rect 21174 14220 21180 14232
rect 21232 14220 21238 14272
rect 24486 14220 24492 14272
rect 24544 14260 24550 14272
rect 26142 14260 26148 14272
rect 24544 14232 26148 14260
rect 24544 14220 24550 14232
rect 26142 14220 26148 14232
rect 26200 14220 26206 14272
rect 27430 14220 27436 14272
rect 27488 14260 27494 14272
rect 29932 14260 29960 14368
rect 30558 14356 30564 14368
rect 30616 14356 30622 14408
rect 30834 14396 30840 14408
rect 30795 14368 30840 14396
rect 30834 14356 30840 14368
rect 30892 14356 30898 14408
rect 31386 14356 31392 14408
rect 31444 14396 31450 14408
rect 31665 14399 31723 14405
rect 31665 14396 31677 14399
rect 31444 14368 31677 14396
rect 31444 14356 31450 14368
rect 31665 14365 31677 14368
rect 31711 14365 31723 14399
rect 31846 14396 31852 14408
rect 31807 14368 31852 14396
rect 31665 14359 31723 14365
rect 31846 14356 31852 14368
rect 31904 14356 31910 14408
rect 32030 14396 32036 14408
rect 31991 14368 32036 14396
rect 32030 14356 32036 14368
rect 32088 14356 32094 14408
rect 32214 14396 32220 14408
rect 32175 14368 32220 14396
rect 32214 14356 32220 14368
rect 32272 14356 32278 14408
rect 32306 14356 32312 14408
rect 32364 14396 32370 14408
rect 33428 14396 33456 14427
rect 47762 14424 47768 14436
rect 47820 14424 47826 14476
rect 32364 14368 33456 14396
rect 32364 14356 32370 14368
rect 30009 14331 30067 14337
rect 30009 14297 30021 14331
rect 30055 14328 30067 14331
rect 30650 14328 30656 14340
rect 30055 14300 30656 14328
rect 30055 14297 30067 14300
rect 30009 14291 30067 14297
rect 30650 14288 30656 14300
rect 30708 14288 30714 14340
rect 27488 14232 29960 14260
rect 27488 14220 27494 14232
rect 30098 14220 30104 14272
rect 30156 14260 30162 14272
rect 32048 14260 32076 14356
rect 33226 14328 33232 14340
rect 33187 14300 33232 14328
rect 33226 14288 33232 14300
rect 33284 14288 33290 14340
rect 46477 14331 46535 14337
rect 46477 14297 46489 14331
rect 46523 14328 46535 14331
rect 46842 14328 46848 14340
rect 46523 14300 46848 14328
rect 46523 14297 46535 14300
rect 46477 14291 46535 14297
rect 46842 14288 46848 14300
rect 46900 14288 46906 14340
rect 48130 14328 48136 14340
rect 48091 14300 48136 14328
rect 48130 14288 48136 14300
rect 48188 14288 48194 14340
rect 30156 14232 32076 14260
rect 32401 14263 32459 14269
rect 30156 14220 30162 14232
rect 32401 14229 32413 14263
rect 32447 14260 32459 14263
rect 32674 14260 32680 14272
rect 32447 14232 32680 14260
rect 32447 14229 32459 14232
rect 32401 14223 32459 14229
rect 32674 14220 32680 14232
rect 32732 14220 32738 14272
rect 1104 14170 48852 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 48852 14170
rect 1104 14096 48852 14118
rect 20162 14056 20168 14068
rect 19628 14028 20168 14056
rect 1762 13920 1768 13932
rect 1723 13892 1768 13920
rect 1762 13880 1768 13892
rect 1820 13880 1826 13932
rect 17034 13880 17040 13932
rect 17092 13920 17098 13932
rect 19628 13929 19656 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 24765 14059 24823 14065
rect 24765 14056 24777 14059
rect 23584 14028 24777 14056
rect 20809 13991 20867 13997
rect 20809 13988 20821 13991
rect 19904 13960 20821 13988
rect 19904 13929 19932 13960
rect 20809 13957 20821 13960
rect 20855 13957 20867 13991
rect 23584 13988 23612 14028
rect 24765 14025 24777 14028
rect 24811 14025 24823 14059
rect 24765 14019 24823 14025
rect 27157 14059 27215 14065
rect 27157 14025 27169 14059
rect 27203 14056 27215 14059
rect 27430 14056 27436 14068
rect 27203 14028 27436 14056
rect 27203 14025 27215 14028
rect 27157 14019 27215 14025
rect 27430 14016 27436 14028
rect 27488 14016 27494 14068
rect 27985 14059 28043 14065
rect 27985 14025 27997 14059
rect 28031 14025 28043 14059
rect 27985 14019 28043 14025
rect 20809 13951 20867 13957
rect 23492 13960 23612 13988
rect 17129 13923 17187 13929
rect 17129 13920 17141 13923
rect 17092 13892 17141 13920
rect 17092 13880 17098 13892
rect 17129 13889 17141 13892
rect 17175 13889 17187 13923
rect 17129 13883 17187 13889
rect 19613 13923 19671 13929
rect 19613 13889 19625 13923
rect 19659 13889 19671 13923
rect 19613 13883 19671 13889
rect 19705 13923 19763 13929
rect 19705 13889 19717 13923
rect 19751 13889 19763 13923
rect 19705 13883 19763 13889
rect 19889 13923 19947 13929
rect 19889 13889 19901 13923
rect 19935 13889 19947 13923
rect 19889 13883 19947 13889
rect 19981 13923 20039 13929
rect 19981 13889 19993 13923
rect 20027 13920 20039 13923
rect 20625 13923 20683 13929
rect 20027 13892 20576 13920
rect 20027 13889 20039 13892
rect 19981 13883 20039 13889
rect 1946 13852 1952 13864
rect 1907 13824 1952 13852
rect 1946 13812 1952 13824
rect 2004 13812 2010 13864
rect 2774 13812 2780 13864
rect 2832 13852 2838 13864
rect 17310 13852 17316 13864
rect 2832 13824 2877 13852
rect 17271 13824 17316 13852
rect 2832 13812 2838 13824
rect 17310 13812 17316 13824
rect 17368 13812 17374 13864
rect 18046 13852 18052 13864
rect 18007 13824 18052 13852
rect 18046 13812 18052 13824
rect 18104 13812 18110 13864
rect 19426 13812 19432 13864
rect 19484 13852 19490 13864
rect 19720 13852 19748 13883
rect 19484 13824 19748 13852
rect 19484 13812 19490 13824
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 20441 13855 20499 13861
rect 20441 13852 20453 13855
rect 20312 13824 20453 13852
rect 20312 13812 20318 13824
rect 20441 13821 20453 13824
rect 20487 13821 20499 13855
rect 20548 13852 20576 13892
rect 20625 13889 20637 13923
rect 20671 13920 20683 13923
rect 20714 13920 20720 13932
rect 20671 13892 20720 13920
rect 20671 13889 20683 13892
rect 20625 13883 20683 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 23492 13929 23520 13960
rect 23842 13948 23848 14000
rect 23900 13988 23906 14000
rect 24397 13991 24455 13997
rect 24397 13988 24409 13991
rect 23900 13960 24409 13988
rect 23900 13948 23906 13960
rect 24397 13957 24409 13960
rect 24443 13957 24455 13991
rect 24397 13951 24455 13957
rect 24486 13948 24492 14000
rect 24544 13988 24550 14000
rect 24597 13991 24655 13997
rect 24597 13988 24609 13991
rect 24544 13960 24609 13988
rect 24544 13948 24550 13960
rect 24597 13957 24609 13960
rect 24643 13957 24655 13991
rect 25501 13991 25559 13997
rect 25501 13988 25513 13991
rect 24597 13951 24655 13957
rect 24688 13960 25513 13988
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 23569 13923 23627 13929
rect 23569 13889 23581 13923
rect 23615 13920 23627 13923
rect 24688 13920 24716 13960
rect 25501 13957 25513 13960
rect 25547 13957 25559 13991
rect 25501 13951 25559 13957
rect 26142 13948 26148 14000
rect 26200 13988 26206 14000
rect 26237 13991 26295 13997
rect 26237 13988 26249 13991
rect 26200 13960 26249 13988
rect 26200 13948 26206 13960
rect 26237 13957 26249 13960
rect 26283 13957 26295 13991
rect 26237 13951 26295 13957
rect 26421 13991 26479 13997
rect 26421 13957 26433 13991
rect 26467 13988 26479 13991
rect 26878 13988 26884 14000
rect 26467 13960 26884 13988
rect 26467 13957 26479 13960
rect 26421 13951 26479 13957
rect 26878 13948 26884 13960
rect 26936 13948 26942 14000
rect 28000 13988 28028 14019
rect 29178 14016 29184 14068
rect 29236 14056 29242 14068
rect 30926 14056 30932 14068
rect 29236 14028 30932 14056
rect 29236 14016 29242 14028
rect 30926 14016 30932 14028
rect 30984 14016 30990 14068
rect 31386 14056 31392 14068
rect 31347 14028 31392 14056
rect 31386 14016 31392 14028
rect 31444 14016 31450 14068
rect 32122 14016 32128 14068
rect 32180 14056 32186 14068
rect 33781 14059 33839 14065
rect 33781 14056 33793 14059
rect 32180 14028 33793 14056
rect 32180 14016 32186 14028
rect 33781 14025 33793 14028
rect 33827 14025 33839 14059
rect 46842 14056 46848 14068
rect 46803 14028 46848 14056
rect 33781 14019 33839 14025
rect 46842 14016 46848 14028
rect 46900 14016 46906 14068
rect 48038 14056 48044 14068
rect 47999 14028 48044 14056
rect 48038 14016 48044 14028
rect 48096 14016 48102 14068
rect 32306 13988 32312 14000
rect 28000 13960 32312 13988
rect 32306 13948 32312 13960
rect 32364 13948 32370 14000
rect 32674 13997 32680 14000
rect 32668 13988 32680 13997
rect 32635 13960 32680 13988
rect 32668 13951 32680 13960
rect 32674 13948 32680 13951
rect 32732 13948 32738 14000
rect 23615 13892 24716 13920
rect 25225 13923 25283 13929
rect 23615 13889 23627 13892
rect 23569 13883 23627 13889
rect 25225 13889 25237 13923
rect 25271 13889 25283 13923
rect 25225 13883 25283 13889
rect 26973 13923 27031 13929
rect 26973 13889 26985 13923
rect 27019 13920 27031 13923
rect 27246 13920 27252 13932
rect 27019 13892 27252 13920
rect 27019 13889 27031 13892
rect 26973 13883 27031 13889
rect 20990 13852 20996 13864
rect 20548 13824 20996 13852
rect 20441 13815 20499 13821
rect 20990 13812 20996 13824
rect 21048 13812 21054 13864
rect 23658 13812 23664 13864
rect 23716 13852 23722 13864
rect 23845 13855 23903 13861
rect 23845 13852 23857 13855
rect 23716 13824 23857 13852
rect 23716 13812 23722 13824
rect 23845 13821 23857 13824
rect 23891 13821 23903 13855
rect 23845 13815 23903 13821
rect 23937 13855 23995 13861
rect 23937 13821 23949 13855
rect 23983 13852 23995 13855
rect 24118 13852 24124 13864
rect 23983 13824 24124 13852
rect 23983 13821 23995 13824
rect 23937 13815 23995 13821
rect 19429 13719 19487 13725
rect 19429 13685 19441 13719
rect 19475 13716 19487 13719
rect 19518 13716 19524 13728
rect 19475 13688 19524 13716
rect 19475 13685 19487 13688
rect 19429 13679 19487 13685
rect 19518 13676 19524 13688
rect 19576 13676 19582 13728
rect 23290 13716 23296 13728
rect 23251 13688 23296 13716
rect 23290 13676 23296 13688
rect 23348 13676 23354 13728
rect 23860 13716 23888 13815
rect 24118 13812 24124 13824
rect 24176 13812 24182 13864
rect 25240 13852 25268 13883
rect 27246 13880 27252 13892
rect 27304 13880 27310 13932
rect 27801 13923 27859 13929
rect 27801 13889 27813 13923
rect 27847 13920 27859 13923
rect 27890 13920 27896 13932
rect 27847 13892 27896 13920
rect 27847 13889 27859 13892
rect 27801 13883 27859 13889
rect 27890 13880 27896 13892
rect 27948 13880 27954 13932
rect 29454 13920 29460 13932
rect 29415 13892 29460 13920
rect 29454 13880 29460 13892
rect 29512 13880 29518 13932
rect 29638 13920 29644 13932
rect 29599 13892 29644 13920
rect 29638 13880 29644 13892
rect 29696 13880 29702 13932
rect 31018 13920 31024 13932
rect 30979 13892 31024 13920
rect 31018 13880 31024 13892
rect 31076 13880 31082 13932
rect 32398 13920 32404 13932
rect 31726 13892 32404 13920
rect 24228 13824 25268 13852
rect 25501 13855 25559 13861
rect 24026 13744 24032 13796
rect 24084 13784 24090 13796
rect 24228 13784 24256 13824
rect 25501 13821 25513 13855
rect 25547 13852 25559 13855
rect 26418 13852 26424 13864
rect 25547 13824 26424 13852
rect 25547 13821 25559 13824
rect 25501 13815 25559 13821
rect 26418 13812 26424 13824
rect 26476 13812 26482 13864
rect 29549 13855 29607 13861
rect 29549 13821 29561 13855
rect 29595 13821 29607 13855
rect 29549 13815 29607 13821
rect 30101 13855 30159 13861
rect 30101 13821 30113 13855
rect 30147 13852 30159 13855
rect 30650 13852 30656 13864
rect 30147 13824 30656 13852
rect 30147 13821 30159 13824
rect 30101 13815 30159 13821
rect 26326 13784 26332 13796
rect 24084 13756 24256 13784
rect 24320 13756 26332 13784
rect 24084 13744 24090 13756
rect 24320 13716 24348 13756
rect 26326 13744 26332 13756
rect 26384 13744 26390 13796
rect 29564 13784 29592 13815
rect 30650 13812 30656 13824
rect 30708 13812 30714 13864
rect 30926 13812 30932 13864
rect 30984 13852 30990 13864
rect 31113 13855 31171 13861
rect 31113 13852 31125 13855
rect 30984 13824 31125 13852
rect 30984 13812 30990 13824
rect 31113 13821 31125 13824
rect 31159 13821 31171 13855
rect 31113 13815 31171 13821
rect 30006 13784 30012 13796
rect 29564 13756 30012 13784
rect 30006 13744 30012 13756
rect 30064 13784 30070 13796
rect 30377 13787 30435 13793
rect 30377 13784 30389 13787
rect 30064 13756 30389 13784
rect 30064 13744 30070 13756
rect 30377 13753 30389 13756
rect 30423 13753 30435 13787
rect 30377 13747 30435 13753
rect 30742 13744 30748 13796
rect 30800 13784 30806 13796
rect 31726 13784 31754 13892
rect 32398 13880 32404 13892
rect 32456 13880 32462 13932
rect 33778 13880 33784 13932
rect 33836 13920 33842 13932
rect 46753 13923 46811 13929
rect 46753 13920 46765 13923
rect 33836 13892 46765 13920
rect 33836 13880 33842 13892
rect 46753 13889 46765 13892
rect 46799 13889 46811 13923
rect 47854 13920 47860 13932
rect 47815 13892 47860 13920
rect 46753 13883 46811 13889
rect 47854 13880 47860 13892
rect 47912 13880 47918 13932
rect 30800 13756 31754 13784
rect 30800 13744 30806 13756
rect 24578 13716 24584 13728
rect 23860 13688 24348 13716
rect 24539 13688 24584 13716
rect 24578 13676 24584 13688
rect 24636 13676 24642 13728
rect 24670 13676 24676 13728
rect 24728 13716 24734 13728
rect 25317 13719 25375 13725
rect 25317 13716 25329 13719
rect 24728 13688 25329 13716
rect 24728 13676 24734 13688
rect 25317 13685 25329 13688
rect 25363 13685 25375 13719
rect 25317 13679 25375 13685
rect 30561 13719 30619 13725
rect 30561 13685 30573 13719
rect 30607 13716 30619 13719
rect 30834 13716 30840 13728
rect 30607 13688 30840 13716
rect 30607 13685 30619 13688
rect 30561 13679 30619 13685
rect 30834 13676 30840 13688
rect 30892 13716 30898 13728
rect 31021 13719 31079 13725
rect 31021 13716 31033 13719
rect 30892 13688 31033 13716
rect 30892 13676 30898 13688
rect 31021 13685 31033 13688
rect 31067 13685 31079 13719
rect 31021 13679 31079 13685
rect 1104 13626 48852 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 48852 13626
rect 1104 13552 48852 13574
rect 1946 13472 1952 13524
rect 2004 13512 2010 13524
rect 2133 13515 2191 13521
rect 2133 13512 2145 13515
rect 2004 13484 2145 13512
rect 2004 13472 2010 13484
rect 2133 13481 2145 13484
rect 2179 13481 2191 13515
rect 17310 13512 17316 13524
rect 17271 13484 17316 13512
rect 2133 13475 2191 13481
rect 17310 13472 17316 13484
rect 17368 13472 17374 13524
rect 21818 13512 21824 13524
rect 17420 13484 21824 13512
rect 1946 13268 1952 13320
rect 2004 13308 2010 13320
rect 2041 13311 2099 13317
rect 2041 13308 2053 13311
rect 2004 13280 2053 13308
rect 2004 13268 2010 13280
rect 2041 13277 2053 13280
rect 2087 13308 2099 13311
rect 2314 13308 2320 13320
rect 2087 13280 2320 13308
rect 2087 13277 2099 13280
rect 2041 13271 2099 13277
rect 2314 13268 2320 13280
rect 2372 13268 2378 13320
rect 7098 13268 7104 13320
rect 7156 13308 7162 13320
rect 16850 13308 16856 13320
rect 7156 13280 16856 13308
rect 7156 13268 7162 13280
rect 16850 13268 16856 13280
rect 16908 13308 16914 13320
rect 17221 13311 17279 13317
rect 17221 13308 17233 13311
rect 16908 13280 17233 13308
rect 16908 13268 16914 13280
rect 17221 13277 17233 13280
rect 17267 13308 17279 13311
rect 17420 13308 17448 13484
rect 21818 13472 21824 13484
rect 21876 13472 21882 13524
rect 23842 13472 23848 13524
rect 23900 13512 23906 13524
rect 24302 13512 24308 13524
rect 23900 13484 24308 13512
rect 23900 13472 23906 13484
rect 24302 13472 24308 13484
rect 24360 13472 24366 13524
rect 27246 13512 27252 13524
rect 24412 13484 27252 13512
rect 24412 13444 24440 13484
rect 27246 13472 27252 13484
rect 27304 13472 27310 13524
rect 29362 13472 29368 13524
rect 29420 13512 29426 13524
rect 29917 13515 29975 13521
rect 29917 13512 29929 13515
rect 29420 13484 29929 13512
rect 29420 13472 29426 13484
rect 29917 13481 29929 13484
rect 29963 13481 29975 13515
rect 29917 13475 29975 13481
rect 30469 13515 30527 13521
rect 30469 13481 30481 13515
rect 30515 13512 30527 13515
rect 31018 13512 31024 13524
rect 30515 13484 31024 13512
rect 30515 13481 30527 13484
rect 30469 13475 30527 13481
rect 31018 13472 31024 13484
rect 31076 13472 31082 13524
rect 23400 13416 24440 13444
rect 19242 13376 19248 13388
rect 19203 13348 19248 13376
rect 19242 13336 19248 13348
rect 19300 13336 19306 13388
rect 19518 13317 19524 13320
rect 19512 13308 19524 13317
rect 17267 13280 17448 13308
rect 19479 13280 19524 13308
rect 17267 13277 17279 13280
rect 17221 13271 17279 13277
rect 19512 13271 19524 13280
rect 19518 13268 19524 13271
rect 19576 13268 19582 13320
rect 21358 13268 21364 13320
rect 21416 13308 21422 13320
rect 22189 13311 22247 13317
rect 22189 13308 22201 13311
rect 21416 13280 22201 13308
rect 21416 13268 21422 13280
rect 22189 13277 22201 13280
rect 22235 13277 22247 13311
rect 22189 13271 22247 13277
rect 22456 13311 22514 13317
rect 22456 13277 22468 13311
rect 22502 13308 22514 13311
rect 23290 13308 23296 13320
rect 22502 13280 23296 13308
rect 22502 13277 22514 13280
rect 22456 13271 22514 13277
rect 23290 13268 23296 13280
rect 23348 13268 23354 13320
rect 20162 13200 20168 13252
rect 20220 13240 20226 13252
rect 23400 13240 23428 13416
rect 25958 13404 25964 13456
rect 26016 13444 26022 13456
rect 26234 13444 26240 13456
rect 26016 13416 26240 13444
rect 26016 13404 26022 13416
rect 26234 13404 26240 13416
rect 26292 13404 26298 13456
rect 29454 13404 29460 13456
rect 29512 13444 29518 13456
rect 30837 13447 30895 13453
rect 30837 13444 30849 13447
rect 29512 13416 30849 13444
rect 29512 13404 29518 13416
rect 30837 13413 30849 13416
rect 30883 13413 30895 13447
rect 30837 13407 30895 13413
rect 23474 13336 23480 13388
rect 23532 13376 23538 13388
rect 24486 13376 24492 13388
rect 23532 13348 24492 13376
rect 23532 13336 23538 13348
rect 24486 13336 24492 13348
rect 24544 13376 24550 13388
rect 24762 13376 24768 13388
rect 24544 13348 24768 13376
rect 24544 13336 24550 13348
rect 24762 13336 24768 13348
rect 24820 13376 24826 13388
rect 25498 13376 25504 13388
rect 24820 13348 25268 13376
rect 25459 13348 25504 13376
rect 24820 13336 24826 13348
rect 24397 13311 24455 13317
rect 24397 13277 24409 13311
rect 24443 13308 24455 13311
rect 24670 13308 24676 13320
rect 24443 13280 24676 13308
rect 24443 13277 24455 13280
rect 24397 13271 24455 13277
rect 24670 13268 24676 13280
rect 24728 13268 24734 13320
rect 25240 13317 25268 13348
rect 25498 13336 25504 13348
rect 25556 13336 25562 13388
rect 27154 13336 27160 13388
rect 27212 13376 27218 13388
rect 28166 13376 28172 13388
rect 27212 13348 28172 13376
rect 27212 13336 27218 13348
rect 28166 13336 28172 13348
rect 28224 13376 28230 13388
rect 30929 13379 30987 13385
rect 30929 13376 30941 13379
rect 28224 13348 30941 13376
rect 28224 13336 28230 13348
rect 30929 13345 30941 13348
rect 30975 13345 30987 13379
rect 32122 13376 32128 13388
rect 32083 13348 32128 13376
rect 30929 13339 30987 13345
rect 32122 13336 32128 13348
rect 32180 13336 32186 13388
rect 32306 13376 32312 13388
rect 32267 13348 32312 13376
rect 32306 13336 32312 13348
rect 32364 13336 32370 13388
rect 25225 13311 25283 13317
rect 25225 13277 25237 13311
rect 25271 13277 25283 13311
rect 25225 13271 25283 13277
rect 25314 13268 25320 13320
rect 25372 13308 25378 13320
rect 26053 13311 26111 13317
rect 25372 13280 25417 13308
rect 25372 13268 25378 13280
rect 26053 13277 26065 13311
rect 26099 13308 26111 13311
rect 27798 13308 27804 13320
rect 26099 13280 27804 13308
rect 26099 13277 26111 13280
rect 26053 13271 26111 13277
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 27890 13268 27896 13320
rect 27948 13308 27954 13320
rect 27948 13280 27993 13308
rect 27948 13268 27954 13280
rect 29270 13268 29276 13320
rect 29328 13308 29334 13320
rect 29733 13311 29791 13317
rect 29733 13308 29745 13311
rect 29328 13280 29745 13308
rect 29328 13268 29334 13280
rect 29733 13277 29745 13280
rect 29779 13277 29791 13311
rect 29733 13271 29791 13277
rect 30009 13311 30067 13317
rect 30009 13277 30021 13311
rect 30055 13277 30067 13311
rect 30650 13308 30656 13320
rect 30563 13280 30656 13308
rect 30009 13271 30067 13277
rect 20220 13212 23428 13240
rect 24581 13243 24639 13249
rect 20220 13200 20226 13212
rect 24581 13209 24593 13243
rect 24627 13209 24639 13243
rect 24581 13203 24639 13209
rect 19150 13132 19156 13184
rect 19208 13172 19214 13184
rect 20254 13172 20260 13184
rect 19208 13144 20260 13172
rect 19208 13132 19214 13144
rect 20254 13132 20260 13144
rect 20312 13172 20318 13184
rect 20625 13175 20683 13181
rect 20625 13172 20637 13175
rect 20312 13144 20637 13172
rect 20312 13132 20318 13144
rect 20625 13141 20637 13144
rect 20671 13172 20683 13175
rect 23382 13172 23388 13184
rect 20671 13144 23388 13172
rect 20671 13141 20683 13144
rect 20625 13135 20683 13141
rect 23382 13132 23388 13144
rect 23440 13132 23446 13184
rect 23569 13175 23627 13181
rect 23569 13141 23581 13175
rect 23615 13172 23627 13175
rect 24118 13172 24124 13184
rect 23615 13144 24124 13172
rect 23615 13141 23627 13144
rect 23569 13135 23627 13141
rect 24118 13132 24124 13144
rect 24176 13132 24182 13184
rect 24596 13172 24624 13203
rect 24946 13172 24952 13184
rect 24596 13144 24952 13172
rect 24946 13132 24952 13144
rect 25004 13132 25010 13184
rect 25501 13175 25559 13181
rect 25501 13141 25513 13175
rect 25547 13172 25559 13175
rect 27246 13172 27252 13184
rect 25547 13144 27252 13172
rect 25547 13141 25559 13144
rect 25501 13135 25559 13141
rect 27246 13132 27252 13144
rect 27304 13132 27310 13184
rect 27890 13132 27896 13184
rect 27948 13172 27954 13184
rect 27985 13175 28043 13181
rect 27985 13172 27997 13175
rect 27948 13144 27997 13172
rect 27948 13132 27954 13144
rect 27985 13141 27997 13144
rect 28031 13141 28043 13175
rect 27985 13135 28043 13141
rect 29549 13175 29607 13181
rect 29549 13141 29561 13175
rect 29595 13172 29607 13175
rect 29638 13172 29644 13184
rect 29595 13144 29644 13172
rect 29595 13141 29607 13144
rect 29549 13135 29607 13141
rect 29638 13132 29644 13144
rect 29696 13132 29702 13184
rect 30024 13172 30052 13271
rect 30650 13268 30656 13280
rect 30708 13268 30714 13320
rect 32033 13311 32091 13317
rect 32033 13277 32045 13311
rect 32079 13308 32091 13311
rect 32214 13308 32220 13320
rect 32079 13280 32220 13308
rect 32079 13277 32091 13280
rect 32033 13271 32091 13277
rect 32214 13268 32220 13280
rect 32272 13268 32278 13320
rect 30668 13240 30696 13268
rect 30668 13212 31708 13240
rect 30558 13172 30564 13184
rect 30024 13144 30564 13172
rect 30558 13132 30564 13144
rect 30616 13172 30622 13184
rect 31110 13172 31116 13184
rect 30616 13144 31116 13172
rect 30616 13132 30622 13144
rect 31110 13132 31116 13144
rect 31168 13132 31174 13184
rect 31680 13181 31708 13212
rect 31665 13175 31723 13181
rect 31665 13141 31677 13175
rect 31711 13141 31723 13175
rect 31665 13135 31723 13141
rect 32306 13132 32312 13184
rect 32364 13172 32370 13184
rect 32766 13172 32772 13184
rect 32364 13144 32772 13172
rect 32364 13132 32370 13144
rect 32766 13132 32772 13144
rect 32824 13132 32830 13184
rect 1104 13082 48852 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 48852 13082
rect 1104 13008 48852 13030
rect 23474 12968 23480 12980
rect 22204 12940 23480 12968
rect 1673 12835 1731 12841
rect 1673 12801 1685 12835
rect 1719 12832 1731 12835
rect 3510 12832 3516 12844
rect 1719 12804 3516 12832
rect 1719 12801 1731 12804
rect 1673 12795 1731 12801
rect 3510 12792 3516 12804
rect 3568 12792 3574 12844
rect 16850 12832 16856 12844
rect 16811 12804 16856 12832
rect 16850 12792 16856 12804
rect 16908 12792 16914 12844
rect 18230 12832 18236 12844
rect 18191 12804 18236 12832
rect 18230 12792 18236 12804
rect 18288 12792 18294 12844
rect 18509 12835 18567 12841
rect 18509 12801 18521 12835
rect 18555 12832 18567 12835
rect 19242 12832 19248 12844
rect 18555 12804 19248 12832
rect 18555 12801 18567 12804
rect 18509 12795 18567 12801
rect 19242 12792 19248 12804
rect 19300 12832 19306 12844
rect 20809 12835 20867 12841
rect 20809 12832 20821 12835
rect 19300 12804 20821 12832
rect 19300 12792 19306 12804
rect 20809 12801 20821 12804
rect 20855 12801 20867 12835
rect 20809 12795 20867 12801
rect 20993 12835 21051 12841
rect 20993 12801 21005 12835
rect 21039 12832 21051 12835
rect 21266 12832 21272 12844
rect 21039 12804 21272 12832
rect 21039 12801 21051 12804
rect 20993 12795 21051 12801
rect 21266 12792 21272 12804
rect 21324 12792 21330 12844
rect 22204 12841 22232 12940
rect 23474 12928 23480 12940
rect 23532 12928 23538 12980
rect 24762 12928 24768 12980
rect 24820 12968 24826 12980
rect 25225 12971 25283 12977
rect 25225 12968 25237 12971
rect 24820 12940 25237 12968
rect 24820 12928 24826 12940
rect 25225 12937 25237 12940
rect 25271 12937 25283 12971
rect 27154 12968 27160 12980
rect 27115 12940 27160 12968
rect 25225 12931 25283 12937
rect 27154 12928 27160 12940
rect 27212 12928 27218 12980
rect 24857 12903 24915 12909
rect 24857 12900 24869 12903
rect 22940 12872 24869 12900
rect 22940 12841 22968 12872
rect 24857 12869 24869 12872
rect 24903 12869 24915 12903
rect 24857 12863 24915 12869
rect 25590 12860 25596 12912
rect 25648 12900 25654 12912
rect 26145 12903 26203 12909
rect 26145 12900 26157 12903
rect 25648 12872 26157 12900
rect 25648 12860 25654 12872
rect 26145 12869 26157 12872
rect 26191 12869 26203 12903
rect 26145 12863 26203 12869
rect 26973 12903 27031 12909
rect 26973 12869 26985 12903
rect 27019 12900 27031 12903
rect 27614 12900 27620 12912
rect 27019 12872 27620 12900
rect 27019 12869 27031 12872
rect 26973 12863 27031 12869
rect 27614 12860 27620 12872
rect 27672 12860 27678 12912
rect 27798 12860 27804 12912
rect 27856 12900 27862 12912
rect 28997 12903 29055 12909
rect 28997 12900 29009 12903
rect 27856 12872 29009 12900
rect 27856 12860 27862 12872
rect 28997 12869 29009 12872
rect 29043 12869 29055 12903
rect 28997 12863 29055 12869
rect 29917 12903 29975 12909
rect 29917 12869 29929 12903
rect 29963 12900 29975 12903
rect 30650 12900 30656 12912
rect 29963 12872 30656 12900
rect 29963 12869 29975 12872
rect 29917 12863 29975 12869
rect 30650 12860 30656 12872
rect 30708 12860 30714 12912
rect 36633 12903 36691 12909
rect 36633 12869 36645 12903
rect 36679 12900 36691 12903
rect 37461 12903 37519 12909
rect 37461 12900 37473 12903
rect 36679 12872 37473 12900
rect 36679 12869 36691 12872
rect 36633 12863 36691 12869
rect 37461 12869 37473 12872
rect 37507 12869 37519 12903
rect 37461 12863 37519 12869
rect 22005 12835 22063 12841
rect 22005 12801 22017 12835
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22189 12835 22247 12841
rect 22189 12801 22201 12835
rect 22235 12801 22247 12835
rect 22189 12795 22247 12801
rect 22833 12835 22891 12841
rect 22833 12801 22845 12835
rect 22879 12801 22891 12835
rect 22833 12795 22891 12801
rect 22925 12835 22983 12841
rect 22925 12801 22937 12835
rect 22971 12801 22983 12835
rect 23198 12832 23204 12844
rect 23159 12804 23204 12832
rect 22925 12795 22983 12801
rect 1394 12764 1400 12776
rect 1355 12736 1400 12764
rect 1394 12724 1400 12736
rect 1452 12724 1458 12776
rect 15838 12724 15844 12776
rect 15896 12764 15902 12776
rect 19521 12767 19579 12773
rect 19521 12764 19533 12767
rect 15896 12736 19533 12764
rect 15896 12724 15902 12736
rect 19521 12733 19533 12736
rect 19567 12733 19579 12767
rect 19521 12727 19579 12733
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20254 12764 20260 12776
rect 19843 12736 20260 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 19536 12696 19564 12727
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20162 12696 20168 12708
rect 19536 12668 20168 12696
rect 20162 12656 20168 12668
rect 20220 12656 20226 12708
rect 22020 12696 22048 12795
rect 22097 12767 22155 12773
rect 22097 12733 22109 12767
rect 22143 12764 22155 12767
rect 22848 12764 22876 12795
rect 23198 12792 23204 12804
rect 23256 12792 23262 12844
rect 23290 12792 23296 12844
rect 23348 12832 23354 12844
rect 24026 12832 24032 12844
rect 23348 12804 24032 12832
rect 23348 12792 23354 12804
rect 24026 12792 24032 12804
rect 24084 12792 24090 12844
rect 24394 12792 24400 12844
rect 24452 12832 24458 12844
rect 25041 12835 25099 12841
rect 25041 12832 25053 12835
rect 24452 12804 25053 12832
rect 24452 12792 24458 12804
rect 25041 12801 25053 12804
rect 25087 12801 25099 12835
rect 25041 12795 25099 12801
rect 25314 12792 25320 12844
rect 25372 12832 25378 12844
rect 25777 12835 25835 12841
rect 25372 12804 25417 12832
rect 25372 12792 25378 12804
rect 25777 12801 25789 12835
rect 25823 12801 25835 12835
rect 25777 12795 25835 12801
rect 25925 12835 25983 12841
rect 25925 12801 25937 12835
rect 25971 12832 25983 12835
rect 26053 12835 26111 12841
rect 25971 12801 26004 12832
rect 25925 12795 26004 12801
rect 26053 12801 26065 12835
rect 26099 12822 26111 12835
rect 26099 12801 26188 12822
rect 26053 12795 26188 12801
rect 22143 12736 22876 12764
rect 23109 12767 23167 12773
rect 22143 12733 22155 12736
rect 22097 12727 22155 12733
rect 23109 12733 23121 12767
rect 23155 12764 23167 12767
rect 23842 12764 23848 12776
rect 23155 12736 23848 12764
rect 23155 12733 23167 12736
rect 23109 12727 23167 12733
rect 23842 12724 23848 12736
rect 23900 12724 23906 12776
rect 24118 12764 24124 12776
rect 24079 12736 24124 12764
rect 24118 12724 24124 12736
rect 24176 12724 24182 12776
rect 24305 12767 24363 12773
rect 24305 12733 24317 12767
rect 24351 12764 24363 12767
rect 24486 12764 24492 12776
rect 24351 12736 24492 12764
rect 24351 12733 24363 12736
rect 24305 12727 24363 12733
rect 24486 12724 24492 12736
rect 24544 12724 24550 12776
rect 23474 12696 23480 12708
rect 22020 12668 23480 12696
rect 23474 12656 23480 12668
rect 23532 12656 23538 12708
rect 16942 12628 16948 12640
rect 16903 12600 16948 12628
rect 16942 12588 16948 12600
rect 17000 12588 17006 12640
rect 20714 12588 20720 12640
rect 20772 12628 20778 12640
rect 21177 12631 21235 12637
rect 21177 12628 21189 12631
rect 20772 12600 21189 12628
rect 20772 12588 20778 12600
rect 21177 12597 21189 12600
rect 21223 12597 21235 12631
rect 22646 12628 22652 12640
rect 22607 12600 22652 12628
rect 21177 12591 21235 12597
rect 22646 12588 22652 12600
rect 22704 12588 22710 12640
rect 23658 12628 23664 12640
rect 23571 12600 23664 12628
rect 23658 12588 23664 12600
rect 23716 12628 23722 12640
rect 24670 12628 24676 12640
rect 23716 12600 24676 12628
rect 23716 12588 23722 12600
rect 24670 12588 24676 12600
rect 24728 12588 24734 12640
rect 25792 12628 25820 12795
rect 25976 12696 26004 12795
rect 26068 12794 26188 12795
rect 26160 12764 26188 12794
rect 26234 12792 26240 12844
rect 26292 12841 26298 12844
rect 26292 12832 26300 12841
rect 26292 12804 26337 12832
rect 26292 12795 26300 12804
rect 26292 12792 26298 12795
rect 27246 12792 27252 12844
rect 27304 12832 27310 12844
rect 29638 12832 29644 12844
rect 27304 12804 27349 12832
rect 29599 12804 29644 12832
rect 27304 12792 27310 12804
rect 29638 12792 29644 12804
rect 29696 12792 29702 12844
rect 29822 12832 29828 12844
rect 29783 12804 29828 12832
rect 29822 12792 29828 12804
rect 29880 12792 29886 12844
rect 30009 12835 30067 12841
rect 30009 12801 30021 12835
rect 30055 12801 30067 12835
rect 30009 12795 30067 12801
rect 26326 12764 26332 12776
rect 26160 12736 26332 12764
rect 26326 12724 26332 12736
rect 26384 12764 26390 12776
rect 26384 12736 28994 12764
rect 26384 12724 26390 12736
rect 26142 12696 26148 12708
rect 25976 12668 26148 12696
rect 26142 12656 26148 12668
rect 26200 12656 26206 12708
rect 26973 12699 27031 12705
rect 26973 12696 26985 12699
rect 26252 12668 26985 12696
rect 26252 12628 26280 12668
rect 26973 12665 26985 12668
rect 27019 12665 27031 12699
rect 28966 12696 28994 12736
rect 29730 12724 29736 12776
rect 29788 12764 29794 12776
rect 30024 12764 30052 12795
rect 30190 12792 30196 12844
rect 30248 12832 30254 12844
rect 36541 12835 36599 12841
rect 36541 12832 36553 12835
rect 30248 12804 36553 12832
rect 30248 12792 30254 12804
rect 36541 12801 36553 12804
rect 36587 12801 36599 12835
rect 36541 12795 36599 12801
rect 29788 12736 30052 12764
rect 29788 12724 29794 12736
rect 29748 12696 29776 12724
rect 30742 12696 30748 12708
rect 28966 12668 29776 12696
rect 30116 12668 30748 12696
rect 26973 12659 27031 12665
rect 26418 12628 26424 12640
rect 25792 12600 26280 12628
rect 26379 12600 26424 12628
rect 26418 12588 26424 12600
rect 26476 12588 26482 12640
rect 26878 12588 26884 12640
rect 26936 12628 26942 12640
rect 27154 12628 27160 12640
rect 26936 12600 27160 12628
rect 26936 12588 26942 12600
rect 27154 12588 27160 12600
rect 27212 12588 27218 12640
rect 29089 12631 29147 12637
rect 29089 12597 29101 12631
rect 29135 12628 29147 12631
rect 30116 12628 30144 12668
rect 30742 12656 30748 12668
rect 30800 12656 30806 12708
rect 36556 12696 36584 12795
rect 36630 12724 36636 12776
rect 36688 12764 36694 12776
rect 37277 12767 37335 12773
rect 37277 12764 37289 12767
rect 36688 12736 37289 12764
rect 36688 12724 36694 12736
rect 37277 12733 37289 12736
rect 37323 12733 37335 12767
rect 37277 12727 37335 12733
rect 39117 12767 39175 12773
rect 39117 12733 39129 12767
rect 39163 12764 39175 12767
rect 46842 12764 46848 12776
rect 39163 12736 46848 12764
rect 39163 12733 39175 12736
rect 39117 12727 39175 12733
rect 46842 12724 46848 12736
rect 46900 12724 46906 12776
rect 37826 12696 37832 12708
rect 36556 12668 37832 12696
rect 37826 12656 37832 12668
rect 37884 12656 37890 12708
rect 29135 12600 30144 12628
rect 30193 12631 30251 12637
rect 29135 12597 29147 12600
rect 29089 12591 29147 12597
rect 30193 12597 30205 12631
rect 30239 12628 30251 12631
rect 30834 12628 30840 12640
rect 30239 12600 30840 12628
rect 30239 12597 30251 12600
rect 30193 12591 30251 12597
rect 30834 12588 30840 12600
rect 30892 12588 30898 12640
rect 1104 12538 48852 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 48852 12538
rect 1104 12464 48852 12486
rect 21177 12427 21235 12433
rect 21177 12393 21189 12427
rect 21223 12424 21235 12427
rect 21266 12424 21272 12436
rect 21223 12396 21272 12424
rect 21223 12393 21235 12396
rect 21177 12387 21235 12393
rect 21266 12384 21272 12396
rect 21324 12384 21330 12436
rect 24670 12424 24676 12436
rect 24631 12396 24676 12424
rect 24670 12384 24676 12396
rect 24728 12384 24734 12436
rect 25133 12427 25191 12433
rect 25133 12393 25145 12427
rect 25179 12424 25191 12427
rect 28074 12424 28080 12436
rect 25179 12396 28080 12424
rect 25179 12393 25191 12396
rect 25133 12387 25191 12393
rect 28074 12384 28080 12396
rect 28132 12384 28138 12436
rect 29549 12427 29607 12433
rect 29549 12393 29561 12427
rect 29595 12424 29607 12427
rect 29822 12424 29828 12436
rect 29595 12396 29828 12424
rect 29595 12393 29607 12396
rect 29549 12387 29607 12393
rect 29822 12384 29828 12396
rect 29880 12384 29886 12436
rect 36446 12384 36452 12436
rect 36504 12424 36510 12436
rect 45554 12424 45560 12436
rect 36504 12396 45560 12424
rect 36504 12384 36510 12396
rect 45554 12384 45560 12396
rect 45612 12384 45618 12436
rect 23753 12359 23811 12365
rect 23753 12325 23765 12359
rect 23799 12356 23811 12359
rect 24578 12356 24584 12368
rect 23799 12328 24584 12356
rect 23799 12325 23811 12328
rect 23753 12319 23811 12325
rect 24578 12316 24584 12328
rect 24636 12316 24642 12368
rect 25038 12356 25044 12368
rect 24688 12328 25044 12356
rect 22646 12248 22652 12300
rect 22704 12288 22710 12300
rect 22925 12291 22983 12297
rect 22925 12288 22937 12291
rect 22704 12260 22937 12288
rect 22704 12248 22710 12260
rect 22925 12257 22937 12260
rect 22971 12257 22983 12291
rect 22925 12251 22983 12257
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12288 23167 12291
rect 24688 12288 24716 12328
rect 25038 12316 25044 12328
rect 25096 12316 25102 12368
rect 27246 12316 27252 12368
rect 27304 12356 27310 12368
rect 27304 12328 30144 12356
rect 27304 12316 27310 12328
rect 23155 12260 24716 12288
rect 24857 12291 24915 12297
rect 23155 12257 23167 12260
rect 23109 12251 23167 12257
rect 24857 12257 24869 12291
rect 24903 12288 24915 12291
rect 25314 12288 25320 12300
rect 24903 12260 25320 12288
rect 24903 12257 24915 12260
rect 24857 12251 24915 12257
rect 25314 12248 25320 12260
rect 25372 12248 25378 12300
rect 27172 12260 29592 12288
rect 18509 12223 18567 12229
rect 18509 12189 18521 12223
rect 18555 12220 18567 12223
rect 19334 12220 19340 12232
rect 18555 12192 19340 12220
rect 18555 12189 18567 12192
rect 18509 12183 18567 12189
rect 19334 12180 19340 12192
rect 19392 12180 19398 12232
rect 19797 12223 19855 12229
rect 19797 12189 19809 12223
rect 19843 12220 19855 12223
rect 21358 12220 21364 12232
rect 19843 12192 21364 12220
rect 19843 12189 19855 12192
rect 19797 12183 19855 12189
rect 18693 12155 18751 12161
rect 18693 12121 18705 12155
rect 18739 12152 18751 12155
rect 19812 12152 19840 12183
rect 21358 12180 21364 12192
rect 21416 12180 21422 12232
rect 23658 12220 23664 12232
rect 23619 12192 23664 12220
rect 23658 12180 23664 12192
rect 23716 12180 23722 12232
rect 23845 12223 23903 12229
rect 23845 12189 23857 12223
rect 23891 12220 23903 12223
rect 24026 12220 24032 12232
rect 23891 12192 24032 12220
rect 23891 12189 23903 12192
rect 23845 12183 23903 12189
rect 24026 12180 24032 12192
rect 24084 12220 24090 12232
rect 24946 12220 24952 12232
rect 24084 12192 24952 12220
rect 24084 12180 24090 12192
rect 24946 12180 24952 12192
rect 25004 12180 25010 12232
rect 26145 12223 26203 12229
rect 26145 12189 26157 12223
rect 26191 12220 26203 12223
rect 27172 12220 27200 12260
rect 26191 12192 27200 12220
rect 26191 12189 26203 12192
rect 26145 12183 26203 12189
rect 27522 12180 27528 12232
rect 27580 12220 27586 12232
rect 28166 12220 28172 12232
rect 27580 12192 28172 12220
rect 27580 12180 27586 12192
rect 28166 12180 28172 12192
rect 28224 12220 28230 12232
rect 28261 12223 28319 12229
rect 28261 12220 28273 12223
rect 28224 12192 28273 12220
rect 28224 12180 28230 12192
rect 28261 12189 28273 12192
rect 28307 12189 28319 12223
rect 29564 12220 29592 12260
rect 29638 12248 29644 12300
rect 29696 12288 29702 12300
rect 29696 12260 29776 12288
rect 29696 12248 29702 12260
rect 29748 12229 29776 12260
rect 29733 12223 29791 12229
rect 29564 12192 29684 12220
rect 28261 12183 28319 12189
rect 18739 12124 19840 12152
rect 20064 12155 20122 12161
rect 18739 12121 18751 12124
rect 18693 12115 18751 12121
rect 20064 12121 20076 12155
rect 20110 12152 20122 12155
rect 20162 12152 20168 12164
rect 20110 12124 20168 12152
rect 20110 12121 20122 12124
rect 20064 12115 20122 12121
rect 20162 12112 20168 12124
rect 20220 12112 20226 12164
rect 24673 12155 24731 12161
rect 24673 12121 24685 12155
rect 24719 12152 24731 12155
rect 24854 12152 24860 12164
rect 24719 12124 24860 12152
rect 24719 12121 24731 12124
rect 24673 12115 24731 12121
rect 24854 12112 24860 12124
rect 24912 12112 24918 12164
rect 26418 12161 26424 12164
rect 26412 12115 26424 12161
rect 26476 12152 26482 12164
rect 28074 12152 28080 12164
rect 26476 12124 26512 12152
rect 28035 12124 28080 12152
rect 26418 12112 26424 12115
rect 26476 12112 26482 12124
rect 28074 12112 28080 12124
rect 28132 12152 28138 12164
rect 29546 12152 29552 12164
rect 28132 12124 29552 12152
rect 28132 12112 28138 12124
rect 29546 12112 29552 12124
rect 29604 12112 29610 12164
rect 29656 12152 29684 12192
rect 29733 12189 29745 12223
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 29822 12180 29828 12232
rect 29880 12220 29886 12232
rect 30006 12220 30012 12232
rect 29880 12192 29925 12220
rect 29967 12192 30012 12220
rect 29880 12180 29886 12192
rect 30006 12180 30012 12192
rect 30064 12180 30070 12232
rect 30116 12229 30144 12328
rect 30101 12223 30159 12229
rect 30101 12189 30113 12223
rect 30147 12189 30159 12223
rect 30101 12183 30159 12189
rect 30742 12152 30748 12164
rect 29656 12124 30748 12152
rect 30742 12112 30748 12124
rect 30800 12112 30806 12164
rect 22094 12044 22100 12096
rect 22152 12084 22158 12096
rect 22465 12087 22523 12093
rect 22465 12084 22477 12087
rect 22152 12056 22477 12084
rect 22152 12044 22158 12056
rect 22465 12053 22477 12056
rect 22511 12053 22523 12087
rect 22830 12084 22836 12096
rect 22791 12056 22836 12084
rect 22465 12047 22523 12053
rect 22830 12044 22836 12056
rect 22888 12044 22894 12096
rect 23382 12044 23388 12096
rect 23440 12084 23446 12096
rect 25590 12084 25596 12096
rect 23440 12056 25596 12084
rect 23440 12044 23446 12056
rect 25590 12044 25596 12056
rect 25648 12084 25654 12096
rect 26050 12084 26056 12096
rect 25648 12056 26056 12084
rect 25648 12044 25654 12056
rect 26050 12044 26056 12056
rect 26108 12044 26114 12096
rect 26142 12044 26148 12096
rect 26200 12084 26206 12096
rect 27525 12087 27583 12093
rect 27525 12084 27537 12087
rect 26200 12056 27537 12084
rect 26200 12044 26206 12056
rect 27525 12053 27537 12056
rect 27571 12053 27583 12087
rect 27525 12047 27583 12053
rect 1104 11994 48852 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 48852 11994
rect 1104 11920 48852 11942
rect 20162 11880 20168 11892
rect 20123 11852 20168 11880
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 20622 11880 20628 11892
rect 20496 11852 20628 11880
rect 20496 11840 20502 11852
rect 20622 11840 20628 11852
rect 20680 11840 20686 11892
rect 20806 11840 20812 11892
rect 20864 11880 20870 11892
rect 21082 11880 21088 11892
rect 20864 11852 21088 11880
rect 20864 11840 20870 11852
rect 21082 11840 21088 11852
rect 21140 11840 21146 11892
rect 23474 11840 23480 11892
rect 23532 11880 23538 11892
rect 23937 11883 23995 11889
rect 23937 11880 23949 11883
rect 23532 11852 23949 11880
rect 23532 11840 23538 11852
rect 23937 11849 23949 11852
rect 23983 11880 23995 11883
rect 25314 11880 25320 11892
rect 23983 11852 25320 11880
rect 23983 11849 23995 11852
rect 23937 11843 23995 11849
rect 25314 11840 25320 11852
rect 25372 11840 25378 11892
rect 26050 11880 26056 11892
rect 26011 11852 26056 11880
rect 26050 11840 26056 11852
rect 26108 11840 26114 11892
rect 26786 11840 26792 11892
rect 26844 11880 26850 11892
rect 27338 11880 27344 11892
rect 26844 11852 27344 11880
rect 26844 11840 26850 11852
rect 27338 11840 27344 11852
rect 27396 11840 27402 11892
rect 27982 11840 27988 11892
rect 28040 11880 28046 11892
rect 28445 11883 28503 11889
rect 28445 11880 28457 11883
rect 28040 11852 28457 11880
rect 28040 11840 28046 11852
rect 28445 11849 28457 11852
rect 28491 11849 28503 11883
rect 29454 11880 29460 11892
rect 29415 11852 29460 11880
rect 28445 11843 28503 11849
rect 29454 11840 29460 11852
rect 29512 11840 29518 11892
rect 16942 11812 16948 11824
rect 16903 11784 16948 11812
rect 16942 11772 16948 11784
rect 17000 11772 17006 11824
rect 20640 11812 20668 11840
rect 19720 11784 20852 11812
rect 2222 11744 2228 11756
rect 2183 11716 2228 11744
rect 2222 11704 2228 11716
rect 2280 11704 2286 11756
rect 2869 11747 2927 11753
rect 2869 11713 2881 11747
rect 2915 11744 2927 11747
rect 11514 11744 11520 11756
rect 2915 11716 11520 11744
rect 2915 11713 2927 11716
rect 2869 11707 2927 11713
rect 11514 11704 11520 11716
rect 11572 11704 11578 11756
rect 19337 11747 19395 11753
rect 19337 11744 19349 11747
rect 19260 11716 19349 11744
rect 16758 11676 16764 11688
rect 16719 11648 16764 11676
rect 16758 11636 16764 11648
rect 16816 11636 16822 11688
rect 18138 11676 18144 11688
rect 18099 11648 18144 11676
rect 18138 11636 18144 11648
rect 18196 11636 18202 11688
rect 19260 11608 19288 11716
rect 19337 11713 19349 11716
rect 19383 11713 19395 11747
rect 19337 11707 19395 11713
rect 19426 11747 19484 11753
rect 19426 11713 19438 11747
rect 19472 11713 19484 11747
rect 19426 11707 19484 11713
rect 19521 11747 19579 11753
rect 19521 11713 19533 11747
rect 19567 11744 19579 11747
rect 19610 11744 19616 11756
rect 19567 11716 19616 11744
rect 19567 11713 19579 11716
rect 19521 11707 19579 11713
rect 19441 11676 19469 11707
rect 19610 11704 19616 11716
rect 19668 11704 19674 11756
rect 19720 11753 19748 11784
rect 19705 11747 19763 11753
rect 19705 11713 19717 11747
rect 19751 11713 19763 11747
rect 19705 11707 19763 11713
rect 20162 11704 20168 11756
rect 20220 11744 20226 11756
rect 20395 11747 20453 11753
rect 20395 11744 20407 11747
rect 20220 11716 20407 11744
rect 20220 11704 20226 11716
rect 20395 11713 20407 11716
rect 20441 11713 20453 11747
rect 20395 11707 20453 11713
rect 20533 11747 20591 11753
rect 20533 11713 20545 11747
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20625 11747 20683 11753
rect 20625 11713 20637 11747
rect 20671 11744 20683 11747
rect 20714 11744 20720 11756
rect 20671 11716 20720 11744
rect 20671 11713 20683 11716
rect 20625 11707 20683 11713
rect 20254 11676 20260 11688
rect 19441 11648 20260 11676
rect 20254 11636 20260 11648
rect 20312 11676 20318 11688
rect 20548 11676 20576 11707
rect 20714 11704 20720 11716
rect 20772 11704 20778 11756
rect 20824 11753 20852 11784
rect 21266 11772 21272 11824
rect 21324 11812 21330 11824
rect 21324 11784 35894 11812
rect 21324 11772 21330 11784
rect 20809 11747 20867 11753
rect 20809 11713 20821 11747
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 22094 11704 22100 11756
rect 22152 11744 22158 11756
rect 23198 11744 23204 11756
rect 22152 11716 22197 11744
rect 22296 11716 23204 11744
rect 22152 11704 22158 11716
rect 20312 11648 20576 11676
rect 20312 11636 20318 11648
rect 19260 11580 19472 11608
rect 1578 11500 1584 11552
rect 1636 11540 1642 11552
rect 2317 11543 2375 11549
rect 2317 11540 2329 11543
rect 1636 11512 2329 11540
rect 1636 11500 1642 11512
rect 2317 11509 2329 11512
rect 2363 11509 2375 11543
rect 2958 11540 2964 11552
rect 2919 11512 2964 11540
rect 2317 11503 2375 11509
rect 2958 11500 2964 11512
rect 3016 11500 3022 11552
rect 19058 11540 19064 11552
rect 19019 11512 19064 11540
rect 19058 11500 19064 11512
rect 19116 11500 19122 11552
rect 19444 11540 19472 11580
rect 20162 11568 20168 11620
rect 20220 11608 20226 11620
rect 22296 11608 22324 11716
rect 23198 11704 23204 11716
rect 23256 11744 23262 11756
rect 24305 11747 24363 11753
rect 24305 11744 24317 11747
rect 23256 11716 24317 11744
rect 23256 11704 23262 11716
rect 24305 11713 24317 11716
rect 24351 11744 24363 11747
rect 25038 11744 25044 11756
rect 24351 11716 25044 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 25038 11704 25044 11716
rect 25096 11704 25102 11756
rect 25774 11704 25780 11756
rect 25832 11744 25838 11756
rect 27062 11744 27068 11756
rect 25832 11716 27068 11744
rect 25832 11704 25838 11716
rect 27062 11704 27068 11716
rect 27120 11704 27126 11756
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 28261 11747 28319 11753
rect 28261 11744 28273 11747
rect 27672 11716 28273 11744
rect 27672 11704 27678 11716
rect 28261 11713 28273 11716
rect 28307 11713 28319 11747
rect 28261 11707 28319 11713
rect 28537 11747 28595 11753
rect 28537 11713 28549 11747
rect 28583 11713 28595 11747
rect 28537 11707 28595 11713
rect 28997 11747 29055 11753
rect 28997 11713 29009 11747
rect 29043 11744 29055 11747
rect 29043 11716 29224 11744
rect 29043 11713 29055 11716
rect 28997 11707 29055 11713
rect 22830 11636 22836 11688
rect 22888 11676 22894 11688
rect 24397 11679 24455 11685
rect 24397 11676 24409 11679
rect 22888 11648 24409 11676
rect 22888 11636 22894 11648
rect 24397 11645 24409 11648
rect 24443 11645 24455 11679
rect 24397 11639 24455 11645
rect 24486 11636 24492 11688
rect 24544 11676 24550 11688
rect 24581 11679 24639 11685
rect 24581 11676 24593 11679
rect 24544 11648 24593 11676
rect 24544 11636 24550 11648
rect 24581 11645 24593 11648
rect 24627 11676 24639 11679
rect 24670 11676 24676 11688
rect 24627 11648 24676 11676
rect 24627 11645 24639 11648
rect 24581 11639 24639 11645
rect 24670 11636 24676 11648
rect 24728 11636 24734 11688
rect 25590 11636 25596 11688
rect 25648 11676 25654 11688
rect 26142 11676 26148 11688
rect 25648 11648 26148 11676
rect 25648 11636 25654 11648
rect 26142 11636 26148 11648
rect 26200 11636 26206 11688
rect 26326 11676 26332 11688
rect 26287 11648 26332 11676
rect 26326 11636 26332 11648
rect 26384 11636 26390 11688
rect 28552 11676 28580 11707
rect 29089 11679 29147 11685
rect 29089 11676 29101 11679
rect 28552 11648 29101 11676
rect 29089 11645 29101 11648
rect 29135 11645 29147 11679
rect 29196 11676 29224 11716
rect 29270 11704 29276 11756
rect 29328 11744 29334 11756
rect 29328 11716 29373 11744
rect 29328 11704 29334 11716
rect 30466 11704 30472 11756
rect 30524 11744 30530 11756
rect 30561 11747 30619 11753
rect 30561 11744 30573 11747
rect 30524 11716 30573 11744
rect 30524 11704 30530 11716
rect 30561 11713 30573 11716
rect 30607 11713 30619 11747
rect 35866 11744 35894 11784
rect 36630 11744 36636 11756
rect 35866 11716 36636 11744
rect 30561 11707 30619 11713
rect 36630 11704 36636 11716
rect 36688 11704 36694 11756
rect 29638 11676 29644 11688
rect 29196 11648 29644 11676
rect 29089 11639 29147 11645
rect 20220 11580 22324 11608
rect 20220 11568 20226 11580
rect 24854 11568 24860 11620
rect 24912 11608 24918 11620
rect 25498 11608 25504 11620
rect 24912 11580 25504 11608
rect 24912 11568 24918 11580
rect 25498 11568 25504 11580
rect 25556 11608 25562 11620
rect 25685 11611 25743 11617
rect 25685 11608 25697 11611
rect 25556 11580 25697 11608
rect 25556 11568 25562 11580
rect 25685 11577 25697 11580
rect 25731 11577 25743 11611
rect 25685 11571 25743 11577
rect 28626 11568 28632 11620
rect 28684 11608 28690 11620
rect 29104 11608 29132 11639
rect 29638 11636 29644 11648
rect 29696 11676 29702 11688
rect 30650 11676 30656 11688
rect 29696 11648 29776 11676
rect 30611 11648 30656 11676
rect 29696 11636 29702 11648
rect 29546 11608 29552 11620
rect 28684 11580 29040 11608
rect 29104 11580 29552 11608
rect 28684 11568 28690 11580
rect 21542 11540 21548 11552
rect 19444 11512 21548 11540
rect 21542 11500 21548 11512
rect 21600 11500 21606 11552
rect 21910 11540 21916 11552
rect 21871 11512 21916 11540
rect 21910 11500 21916 11512
rect 21968 11500 21974 11552
rect 28261 11543 28319 11549
rect 28261 11509 28273 11543
rect 28307 11540 28319 11543
rect 28902 11540 28908 11552
rect 28307 11512 28908 11540
rect 28307 11509 28319 11512
rect 28261 11503 28319 11509
rect 28902 11500 28908 11512
rect 28960 11500 28966 11552
rect 29012 11549 29040 11580
rect 29546 11568 29552 11580
rect 29604 11568 29610 11620
rect 28997 11543 29055 11549
rect 28997 11509 29009 11543
rect 29043 11509 29055 11543
rect 29748 11540 29776 11648
rect 30650 11636 30656 11648
rect 30708 11636 30714 11688
rect 30745 11679 30803 11685
rect 30745 11645 30757 11679
rect 30791 11676 30803 11679
rect 32490 11676 32496 11688
rect 30791 11648 32496 11676
rect 30791 11645 30803 11648
rect 30745 11639 30803 11645
rect 30098 11568 30104 11620
rect 30156 11608 30162 11620
rect 30760 11608 30788 11639
rect 32490 11636 32496 11648
rect 32548 11636 32554 11688
rect 30156 11580 30788 11608
rect 30156 11568 30162 11580
rect 30193 11543 30251 11549
rect 30193 11540 30205 11543
rect 29748 11512 30205 11540
rect 28997 11503 29055 11509
rect 30193 11509 30205 11512
rect 30239 11509 30251 11543
rect 30193 11503 30251 11509
rect 46290 11500 46296 11552
rect 46348 11540 46354 11552
rect 47765 11543 47823 11549
rect 47765 11540 47777 11543
rect 46348 11512 47777 11540
rect 46348 11500 46354 11512
rect 47765 11509 47777 11512
rect 47811 11509 47823 11543
rect 47765 11503 47823 11509
rect 1104 11450 48852 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 48852 11450
rect 1104 11376 48852 11398
rect 16758 11296 16764 11348
rect 16816 11336 16822 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 16816 11308 18705 11336
rect 16816 11296 16822 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 19610 11336 19616 11348
rect 19571 11308 19616 11336
rect 18693 11299 18751 11305
rect 1581 11203 1639 11209
rect 1581 11169 1593 11203
rect 1627 11200 1639 11203
rect 2958 11200 2964 11212
rect 1627 11172 2964 11200
rect 1627 11169 1639 11172
rect 1581 11163 1639 11169
rect 2958 11160 2964 11172
rect 3016 11160 3022 11212
rect 3050 11160 3056 11212
rect 3108 11200 3114 11212
rect 18708 11200 18736 11299
rect 19610 11296 19616 11308
rect 19668 11296 19674 11348
rect 22741 11339 22799 11345
rect 22741 11305 22753 11339
rect 22787 11336 22799 11339
rect 22830 11336 22836 11348
rect 22787 11308 22836 11336
rect 22787 11305 22799 11308
rect 22741 11299 22799 11305
rect 22830 11296 22836 11308
rect 22888 11296 22894 11348
rect 24857 11339 24915 11345
rect 24857 11305 24869 11339
rect 24903 11336 24915 11339
rect 25590 11336 25596 11348
rect 24903 11308 25596 11336
rect 24903 11305 24915 11308
rect 24857 11299 24915 11305
rect 25590 11296 25596 11308
rect 25648 11296 25654 11348
rect 25682 11296 25688 11348
rect 25740 11336 25746 11348
rect 25869 11339 25927 11345
rect 25869 11336 25881 11339
rect 25740 11308 25881 11336
rect 25740 11296 25746 11308
rect 25869 11305 25881 11308
rect 25915 11305 25927 11339
rect 25869 11299 25927 11305
rect 26234 11296 26240 11348
rect 26292 11336 26298 11348
rect 27338 11336 27344 11348
rect 26292 11308 27344 11336
rect 26292 11296 26298 11308
rect 27338 11296 27344 11308
rect 27396 11336 27402 11348
rect 27801 11339 27859 11345
rect 27801 11336 27813 11339
rect 27396 11308 27813 11336
rect 27396 11296 27402 11308
rect 27801 11305 27813 11308
rect 27847 11336 27859 11339
rect 28813 11339 28871 11345
rect 28813 11336 28825 11339
rect 27847 11308 28825 11336
rect 27847 11305 27859 11308
rect 27801 11299 27859 11305
rect 28813 11305 28825 11308
rect 28859 11336 28871 11339
rect 29270 11336 29276 11348
rect 28859 11308 29276 11336
rect 28859 11305 28871 11308
rect 28813 11299 28871 11305
rect 29270 11296 29276 11308
rect 29328 11296 29334 11348
rect 30650 11296 30656 11348
rect 30708 11336 30714 11348
rect 32125 11339 32183 11345
rect 32125 11336 32137 11339
rect 30708 11308 32137 11336
rect 30708 11296 30714 11308
rect 32125 11305 32137 11308
rect 32171 11305 32183 11339
rect 32125 11299 32183 11305
rect 22848 11200 22876 11296
rect 25041 11271 25099 11277
rect 25041 11237 25053 11271
rect 25087 11237 25099 11271
rect 25041 11231 25099 11237
rect 24673 11203 24731 11209
rect 24673 11200 24685 11203
rect 3108 11172 3153 11200
rect 18708 11172 19472 11200
rect 22848 11172 24685 11200
rect 3108 11160 3114 11172
rect 1397 11135 1455 11141
rect 1397 11101 1409 11135
rect 1443 11101 1455 11135
rect 17310 11132 17316 11144
rect 17271 11104 17316 11132
rect 1397 11095 1455 11101
rect 1412 11064 1440 11095
rect 17310 11092 17316 11104
rect 17368 11092 17374 11144
rect 17580 11135 17638 11141
rect 17580 11101 17592 11135
rect 17626 11132 17638 11135
rect 19058 11132 19064 11144
rect 17626 11104 19064 11132
rect 17626 11101 17638 11104
rect 17580 11095 17638 11101
rect 19058 11092 19064 11104
rect 19116 11092 19122 11144
rect 19242 11132 19248 11144
rect 19203 11104 19248 11132
rect 19242 11092 19248 11104
rect 19300 11092 19306 11144
rect 19444 11141 19472 11172
rect 24673 11169 24685 11172
rect 24719 11169 24731 11203
rect 24673 11163 24731 11169
rect 19429 11135 19487 11141
rect 19429 11101 19441 11135
rect 19475 11101 19487 11135
rect 19429 11095 19487 11101
rect 21082 11092 21088 11144
rect 21140 11132 21146 11144
rect 21358 11132 21364 11144
rect 21140 11104 21364 11132
rect 21140 11092 21146 11104
rect 21358 11092 21364 11104
rect 21416 11092 21422 11144
rect 21628 11135 21686 11141
rect 21628 11101 21640 11135
rect 21674 11132 21686 11135
rect 21910 11132 21916 11144
rect 21674 11104 21916 11132
rect 21674 11101 21686 11104
rect 21628 11095 21686 11101
rect 21910 11092 21916 11104
rect 21968 11092 21974 11144
rect 24118 11092 24124 11144
rect 24176 11132 24182 11144
rect 24857 11135 24915 11141
rect 24857 11132 24869 11135
rect 24176 11104 24869 11132
rect 24176 11092 24182 11104
rect 24857 11101 24869 11104
rect 24903 11101 24915 11135
rect 25056 11132 25084 11231
rect 27154 11228 27160 11280
rect 27212 11268 27218 11280
rect 27522 11268 27528 11280
rect 27212 11240 27528 11268
rect 27212 11228 27218 11240
rect 27522 11228 27528 11240
rect 27580 11268 27586 11280
rect 27580 11240 28948 11268
rect 27580 11228 27586 11240
rect 26326 11160 26332 11212
rect 26384 11200 26390 11212
rect 26384 11172 28856 11200
rect 26384 11160 26390 11172
rect 25501 11135 25559 11141
rect 25501 11132 25513 11135
rect 25056 11104 25513 11132
rect 24857 11095 24915 11101
rect 25501 11101 25513 11104
rect 25547 11101 25559 11135
rect 27614 11132 27620 11144
rect 27575 11104 27620 11132
rect 25501 11095 25559 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 27801 11135 27859 11141
rect 27801 11101 27813 11135
rect 27847 11132 27859 11135
rect 28074 11132 28080 11144
rect 27847 11104 28080 11132
rect 27847 11101 27859 11104
rect 27801 11095 27859 11101
rect 28074 11092 28080 11104
rect 28132 11092 28138 11144
rect 28626 11132 28632 11144
rect 28539 11104 28632 11132
rect 28626 11092 28632 11104
rect 28684 11092 28690 11144
rect 2866 11064 2872 11076
rect 1412 11036 2872 11064
rect 2866 11024 2872 11036
rect 2924 11024 2930 11076
rect 19518 11024 19524 11076
rect 19576 11064 19582 11076
rect 20438 11064 20444 11076
rect 19576 11036 20444 11064
rect 19576 11024 19582 11036
rect 20438 11024 20444 11036
rect 20496 11024 20502 11076
rect 24394 11064 24400 11076
rect 24355 11036 24400 11064
rect 24394 11024 24400 11036
rect 24452 11024 24458 11076
rect 25685 11067 25743 11073
rect 25685 11033 25697 11067
rect 25731 11064 25743 11067
rect 27522 11064 27528 11076
rect 25731 11036 27528 11064
rect 25731 11033 25743 11036
rect 25685 11027 25743 11033
rect 27522 11024 27528 11036
rect 27580 11024 27586 11076
rect 27632 11064 27660 11092
rect 28644 11064 28672 11092
rect 27632 11036 28672 11064
rect 28828 11064 28856 11172
rect 28920 11141 28948 11240
rect 30098 11200 30104 11212
rect 29748 11172 30104 11200
rect 28905 11135 28963 11141
rect 28905 11101 28917 11135
rect 28951 11101 28963 11135
rect 28905 11095 28963 11101
rect 29748 11064 29776 11172
rect 30098 11160 30104 11172
rect 30156 11160 30162 11212
rect 30742 11200 30748 11212
rect 30703 11172 30748 11200
rect 30742 11160 30748 11172
rect 30800 11160 30806 11212
rect 46290 11200 46296 11212
rect 46251 11172 46296 11200
rect 46290 11160 46296 11172
rect 46348 11160 46354 11212
rect 29914 11132 29920 11144
rect 29875 11104 29920 11132
rect 29914 11092 29920 11104
rect 29972 11132 29978 11144
rect 30282 11132 30288 11144
rect 29972 11104 30288 11132
rect 29972 11092 29978 11104
rect 30282 11092 30288 11104
rect 30340 11092 30346 11144
rect 30834 11092 30840 11144
rect 30892 11132 30898 11144
rect 31001 11135 31059 11141
rect 31001 11132 31013 11135
rect 30892 11104 31013 11132
rect 30892 11092 30898 11104
rect 31001 11101 31013 11104
rect 31047 11101 31059 11135
rect 31001 11095 31059 11101
rect 28828 11036 29776 11064
rect 46477 11067 46535 11073
rect 46477 11033 46489 11067
rect 46523 11064 46535 11067
rect 46934 11064 46940 11076
rect 46523 11036 46940 11064
rect 46523 11033 46535 11036
rect 46477 11027 46535 11033
rect 46934 11024 46940 11036
rect 46992 11024 46998 11076
rect 48130 11064 48136 11076
rect 48091 11036 48136 11064
rect 48130 11024 48136 11036
rect 48188 11024 48194 11076
rect 19978 10956 19984 11008
rect 20036 10996 20042 11008
rect 21266 10996 21272 11008
rect 20036 10968 21272 10996
rect 20036 10956 20042 10968
rect 21266 10956 21272 10968
rect 21324 10956 21330 11008
rect 27982 10996 27988 11008
rect 27943 10968 27988 10996
rect 27982 10956 27988 10968
rect 28040 10956 28046 11008
rect 28442 10996 28448 11008
rect 28403 10968 28448 10996
rect 28442 10956 28448 10968
rect 28500 10956 28506 11008
rect 29546 10996 29552 11008
rect 29507 10968 29552 10996
rect 29546 10956 29552 10968
rect 29604 10956 29610 11008
rect 30006 10996 30012 11008
rect 29967 10968 30012 10996
rect 30006 10956 30012 10968
rect 30064 10956 30070 11008
rect 1104 10906 48852 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 48852 10906
rect 1104 10832 48852 10854
rect 27522 10752 27528 10804
rect 27580 10792 27586 10804
rect 29273 10795 29331 10801
rect 29273 10792 29285 10795
rect 27580 10764 29285 10792
rect 27580 10752 27586 10764
rect 29273 10761 29285 10764
rect 29319 10761 29331 10795
rect 29273 10755 29331 10761
rect 29362 10752 29368 10804
rect 29420 10792 29426 10804
rect 31113 10795 31171 10801
rect 31113 10792 31125 10795
rect 29420 10764 31125 10792
rect 29420 10752 29426 10764
rect 31113 10761 31125 10764
rect 31159 10761 31171 10795
rect 46934 10792 46940 10804
rect 46895 10764 46940 10792
rect 31113 10755 31171 10761
rect 46934 10752 46940 10764
rect 46992 10752 46998 10804
rect 20254 10724 20260 10736
rect 19441 10696 20260 10724
rect 19441 10668 19469 10696
rect 20254 10684 20260 10696
rect 20312 10684 20318 10736
rect 27154 10724 27160 10736
rect 26160 10696 27160 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 1673 10659 1731 10665
rect 1673 10625 1685 10659
rect 1719 10656 1731 10659
rect 14550 10656 14556 10668
rect 1719 10628 14556 10656
rect 1719 10625 1731 10628
rect 1673 10619 1731 10625
rect 14550 10616 14556 10628
rect 14608 10616 14614 10668
rect 19150 10616 19156 10668
rect 19208 10656 19214 10668
rect 19291 10659 19349 10665
rect 19291 10656 19303 10659
rect 19208 10628 19303 10656
rect 19208 10616 19214 10628
rect 19291 10625 19303 10628
rect 19337 10625 19349 10659
rect 19291 10619 19349 10625
rect 19426 10662 19484 10668
rect 19426 10628 19438 10662
rect 19472 10628 19484 10662
rect 19426 10622 19484 10628
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10656 19579 10659
rect 19610 10656 19616 10668
rect 19567 10628 19616 10656
rect 19567 10625 19579 10628
rect 19521 10619 19579 10625
rect 19610 10616 19616 10628
rect 19668 10616 19674 10668
rect 19705 10659 19763 10665
rect 19705 10625 19717 10659
rect 19751 10656 19763 10659
rect 20622 10656 20628 10668
rect 19751 10628 20628 10656
rect 19751 10625 19763 10628
rect 19705 10619 19763 10625
rect 20622 10616 20628 10628
rect 20680 10616 20686 10668
rect 24026 10656 24032 10668
rect 23987 10628 24032 10656
rect 24026 10616 24032 10628
rect 24084 10616 24090 10668
rect 26160 10665 26188 10696
rect 27154 10684 27160 10696
rect 27212 10724 27218 10736
rect 27706 10724 27712 10736
rect 27212 10696 27305 10724
rect 27540 10696 27712 10724
rect 27212 10684 27218 10696
rect 26145 10659 26203 10665
rect 26145 10625 26157 10659
rect 26191 10625 26203 10659
rect 26145 10619 26203 10625
rect 26234 10616 26240 10668
rect 26292 10656 26298 10668
rect 26973 10659 27031 10665
rect 26292 10628 26337 10656
rect 26292 10616 26298 10628
rect 26973 10625 26985 10659
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 27249 10659 27307 10665
rect 27249 10625 27261 10659
rect 27295 10656 27307 10659
rect 27338 10656 27344 10668
rect 27295 10628 27344 10656
rect 27295 10625 27307 10628
rect 27249 10619 27307 10625
rect 2866 10588 2872 10600
rect 2827 10560 2872 10588
rect 2866 10548 2872 10560
rect 2924 10548 2930 10600
rect 23106 10548 23112 10600
rect 23164 10588 23170 10600
rect 24489 10591 24547 10597
rect 24489 10588 24501 10591
rect 23164 10560 24501 10588
rect 23164 10548 23170 10560
rect 24489 10557 24501 10560
rect 24535 10557 24547 10591
rect 24489 10551 24547 10557
rect 26326 10548 26332 10600
rect 26384 10548 26390 10600
rect 26421 10591 26479 10597
rect 26421 10557 26433 10591
rect 26467 10557 26479 10591
rect 26988 10588 27016 10619
rect 27338 10616 27344 10628
rect 27396 10616 27402 10668
rect 26988 10580 27476 10588
rect 27540 10580 27568 10696
rect 27706 10684 27712 10696
rect 27764 10724 27770 10736
rect 28902 10724 28908 10736
rect 27764 10696 28908 10724
rect 27764 10684 27770 10696
rect 28902 10684 28908 10696
rect 28960 10684 28966 10736
rect 29012 10696 29408 10724
rect 28813 10659 28871 10665
rect 28813 10625 28825 10659
rect 28859 10656 28871 10659
rect 29012 10656 29040 10696
rect 29270 10666 29276 10668
rect 29104 10665 29276 10666
rect 28859 10628 29040 10656
rect 29082 10659 29276 10665
rect 28859 10625 28871 10628
rect 28813 10619 28871 10625
rect 29082 10625 29094 10659
rect 29128 10638 29276 10659
rect 29128 10625 29140 10638
rect 29082 10619 29140 10625
rect 29270 10616 29276 10638
rect 29328 10616 29334 10668
rect 29380 10656 29408 10696
rect 29454 10684 29460 10736
rect 29512 10724 29518 10736
rect 29512 10696 29960 10724
rect 29512 10684 29518 10696
rect 29730 10656 29736 10668
rect 29380 10628 29592 10656
rect 29691 10628 29736 10656
rect 26988 10560 27568 10580
rect 26421 10551 26479 10557
rect 27448 10552 27568 10560
rect 28997 10591 29055 10597
rect 28997 10557 29009 10591
rect 29043 10588 29055 10591
rect 29564 10588 29592 10628
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 29932 10665 29960 10696
rect 29917 10659 29975 10665
rect 29917 10625 29929 10659
rect 29963 10625 29975 10659
rect 30282 10656 30288 10668
rect 30243 10628 30288 10656
rect 29917 10619 29975 10625
rect 30282 10616 30288 10628
rect 30340 10616 30346 10668
rect 30558 10616 30564 10668
rect 30616 10656 30622 10668
rect 30926 10656 30932 10668
rect 30616 10628 30932 10656
rect 30616 10616 30622 10628
rect 30926 10616 30932 10628
rect 30984 10656 30990 10668
rect 31021 10659 31079 10665
rect 31021 10656 31033 10659
rect 30984 10628 31033 10656
rect 30984 10616 30990 10628
rect 31021 10625 31033 10628
rect 31067 10625 31079 10659
rect 46842 10656 46848 10668
rect 46803 10628 46848 10656
rect 31021 10619 31079 10625
rect 46842 10616 46848 10628
rect 46900 10616 46906 10668
rect 47762 10656 47768 10668
rect 47723 10628 47768 10656
rect 47762 10616 47768 10628
rect 47820 10616 47826 10668
rect 30006 10588 30012 10600
rect 29043 10560 29500 10588
rect 29564 10560 30012 10588
rect 29043 10557 29055 10560
rect 28997 10551 29055 10557
rect 23474 10480 23480 10532
rect 23532 10520 23538 10532
rect 24578 10520 24584 10532
rect 23532 10492 24584 10520
rect 23532 10480 23538 10492
rect 24578 10480 24584 10492
rect 24636 10480 24642 10532
rect 26344 10520 26372 10548
rect 26160 10492 26372 10520
rect 26436 10520 26464 10551
rect 26973 10523 27031 10529
rect 26973 10520 26985 10523
rect 26436 10492 26985 10520
rect 3510 10452 3516 10464
rect 3471 10424 3516 10452
rect 3510 10412 3516 10424
rect 3568 10412 3574 10464
rect 19058 10452 19064 10464
rect 19019 10424 19064 10452
rect 19058 10412 19064 10424
rect 19116 10412 19122 10464
rect 24305 10455 24363 10461
rect 24305 10421 24317 10455
rect 24351 10452 24363 10455
rect 26160 10452 26188 10492
rect 26973 10489 26985 10492
rect 27019 10489 27031 10523
rect 26973 10483 27031 10489
rect 27062 10480 27068 10532
rect 27120 10520 27126 10532
rect 29472 10520 29500 10560
rect 30006 10548 30012 10560
rect 30064 10548 30070 10600
rect 30098 10548 30104 10600
rect 30156 10588 30162 10600
rect 30156 10560 30201 10588
rect 30156 10548 30162 10560
rect 30650 10520 30656 10532
rect 27120 10492 28948 10520
rect 29472 10492 30656 10520
rect 27120 10480 27126 10492
rect 26326 10452 26332 10464
rect 24351 10424 26188 10452
rect 26287 10424 26332 10452
rect 24351 10421 24363 10424
rect 24305 10415 24363 10421
rect 26326 10412 26332 10424
rect 26384 10412 26390 10464
rect 26510 10412 26516 10464
rect 26568 10452 26574 10464
rect 27338 10452 27344 10464
rect 26568 10424 27344 10452
rect 26568 10412 26574 10424
rect 27338 10412 27344 10424
rect 27396 10452 27402 10464
rect 28813 10455 28871 10461
rect 28813 10452 28825 10455
rect 27396 10424 28825 10452
rect 27396 10412 27402 10424
rect 28813 10421 28825 10424
rect 28859 10421 28871 10455
rect 28920 10452 28948 10492
rect 30650 10480 30656 10492
rect 30708 10480 30714 10532
rect 30926 10480 30932 10532
rect 30984 10520 30990 10532
rect 47949 10523 48007 10529
rect 47949 10520 47961 10523
rect 30984 10492 47961 10520
rect 30984 10480 30990 10492
rect 47949 10489 47961 10492
rect 47995 10489 48007 10523
rect 47949 10483 48007 10489
rect 29362 10452 29368 10464
rect 28920 10424 29368 10452
rect 28813 10415 28871 10421
rect 29362 10412 29368 10424
rect 29420 10412 29426 10464
rect 30469 10455 30527 10461
rect 30469 10421 30481 10455
rect 30515 10452 30527 10455
rect 30834 10452 30840 10464
rect 30515 10424 30840 10452
rect 30515 10421 30527 10424
rect 30469 10415 30527 10421
rect 30834 10412 30840 10424
rect 30892 10412 30898 10464
rect 1104 10362 48852 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 48852 10362
rect 1104 10288 48852 10310
rect 19610 10248 19616 10260
rect 19571 10220 19616 10248
rect 19610 10208 19616 10220
rect 19668 10208 19674 10260
rect 21542 10208 21548 10260
rect 21600 10248 21606 10260
rect 23474 10248 23480 10260
rect 21600 10220 22094 10248
rect 21600 10208 21606 10220
rect 20622 10140 20628 10192
rect 20680 10180 20686 10192
rect 20680 10152 20944 10180
rect 20680 10140 20686 10152
rect 1397 10115 1455 10121
rect 1397 10081 1409 10115
rect 1443 10112 1455 10115
rect 3510 10112 3516 10124
rect 1443 10084 3516 10112
rect 1443 10081 1455 10084
rect 1397 10075 1455 10081
rect 3510 10072 3516 10084
rect 3568 10072 3574 10124
rect 20254 10072 20260 10124
rect 20312 10112 20318 10124
rect 20312 10084 20668 10112
rect 20312 10072 20318 10084
rect 19242 10044 19248 10056
rect 19203 10016 19248 10044
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 20640 10053 20668 10084
rect 20533 10047 20591 10053
rect 20533 10013 20545 10047
rect 20579 10013 20591 10047
rect 20533 10007 20591 10013
rect 20625 10047 20683 10053
rect 20625 10013 20637 10047
rect 20671 10013 20683 10047
rect 20625 10007 20683 10013
rect 1578 9976 1584 9988
rect 1539 9948 1584 9976
rect 1578 9936 1584 9948
rect 1636 9936 1642 9988
rect 3234 9976 3240 9988
rect 3195 9948 3240 9976
rect 3234 9936 3240 9948
rect 3292 9936 3298 9988
rect 19334 9936 19340 9988
rect 19392 9976 19398 9988
rect 19429 9979 19487 9985
rect 19429 9976 19441 9979
rect 19392 9948 19441 9976
rect 19392 9936 19398 9948
rect 19429 9945 19441 9948
rect 19475 9945 19487 9979
rect 20548 9976 20576 10007
rect 20714 10004 20720 10056
rect 20772 10044 20778 10056
rect 20916 10053 20944 10152
rect 22066 10112 22094 10220
rect 23308 10220 23480 10248
rect 22066 10084 23060 10112
rect 20901 10047 20959 10053
rect 20772 10016 20817 10044
rect 20772 10004 20778 10016
rect 20901 10013 20913 10047
rect 20947 10013 20959 10047
rect 20901 10007 20959 10013
rect 23032 9976 23060 10084
rect 23106 10004 23112 10056
rect 23164 10044 23170 10056
rect 23308 10053 23336 10220
rect 23474 10208 23480 10220
rect 23532 10208 23538 10260
rect 24026 10208 24032 10260
rect 24084 10248 24090 10260
rect 24397 10251 24455 10257
rect 24397 10248 24409 10251
rect 24084 10220 24409 10248
rect 24084 10208 24090 10220
rect 24397 10217 24409 10220
rect 24443 10217 24455 10251
rect 24397 10211 24455 10217
rect 26053 10251 26111 10257
rect 26053 10217 26065 10251
rect 26099 10248 26111 10251
rect 26234 10248 26240 10260
rect 26099 10220 26240 10248
rect 26099 10217 26111 10220
rect 26053 10211 26111 10217
rect 26234 10208 26240 10220
rect 26292 10208 26298 10260
rect 26418 10208 26424 10260
rect 26476 10248 26482 10260
rect 28445 10251 28503 10257
rect 28445 10248 28457 10251
rect 26476 10220 28457 10248
rect 26476 10208 26482 10220
rect 28445 10217 28457 10220
rect 28491 10248 28503 10251
rect 28491 10220 29040 10248
rect 28491 10217 28503 10220
rect 28445 10211 28503 10217
rect 24670 10140 24676 10192
rect 24728 10180 24734 10192
rect 27890 10180 27896 10192
rect 24728 10152 27896 10180
rect 24728 10140 24734 10152
rect 23394 10115 23452 10121
rect 23394 10081 23406 10115
rect 23440 10112 23452 10115
rect 24394 10112 24400 10124
rect 23440 10084 24400 10112
rect 23440 10081 23452 10084
rect 23394 10075 23452 10081
rect 24394 10072 24400 10084
rect 24452 10112 24458 10124
rect 25056 10121 25084 10152
rect 24857 10115 24915 10121
rect 24857 10112 24869 10115
rect 24452 10084 24869 10112
rect 24452 10072 24458 10084
rect 24857 10081 24869 10084
rect 24903 10081 24915 10115
rect 24857 10075 24915 10081
rect 25041 10115 25099 10121
rect 25041 10081 25053 10115
rect 25087 10081 25099 10115
rect 26510 10112 26516 10124
rect 26471 10084 26516 10112
rect 25041 10075 25099 10081
rect 26510 10072 26516 10084
rect 26568 10072 26574 10124
rect 26712 10121 26740 10152
rect 27890 10140 27896 10152
rect 27948 10180 27954 10192
rect 28534 10180 28540 10192
rect 27948 10152 28540 10180
rect 27948 10140 27954 10152
rect 28534 10140 28540 10152
rect 28592 10140 28598 10192
rect 29012 10180 29040 10220
rect 29822 10208 29828 10260
rect 29880 10248 29886 10260
rect 29917 10251 29975 10257
rect 29917 10248 29929 10251
rect 29880 10220 29929 10248
rect 29880 10208 29886 10220
rect 29917 10217 29929 10220
rect 29963 10217 29975 10251
rect 29917 10211 29975 10217
rect 30006 10208 30012 10260
rect 30064 10248 30070 10260
rect 31941 10251 31999 10257
rect 31941 10248 31953 10251
rect 30064 10220 31953 10248
rect 30064 10208 30070 10220
rect 31941 10217 31953 10220
rect 31987 10217 31999 10251
rect 31941 10211 31999 10217
rect 30558 10180 30564 10192
rect 29012 10152 30564 10180
rect 30558 10140 30564 10152
rect 30616 10140 30622 10192
rect 26697 10115 26755 10121
rect 26697 10081 26709 10115
rect 26743 10081 26755 10115
rect 26697 10075 26755 10081
rect 28442 10072 28448 10124
rect 28500 10112 28506 10124
rect 28629 10115 28687 10121
rect 28629 10112 28641 10115
rect 28500 10084 28641 10112
rect 28500 10072 28506 10084
rect 28629 10081 28641 10084
rect 28675 10081 28687 10115
rect 28629 10075 28687 10081
rect 29380 10084 29868 10112
rect 23293 10047 23351 10053
rect 23164 10016 23209 10044
rect 23164 10004 23170 10016
rect 23293 10013 23305 10047
rect 23339 10013 23351 10047
rect 23474 10044 23480 10056
rect 23435 10016 23480 10044
rect 23293 10007 23351 10013
rect 23474 10004 23480 10016
rect 23532 10004 23538 10056
rect 23661 10047 23719 10053
rect 23661 10042 23673 10047
rect 23584 10014 23673 10042
rect 23584 9976 23612 10014
rect 23661 10013 23673 10014
rect 23707 10044 23719 10047
rect 24765 10047 24823 10053
rect 24765 10044 24777 10047
rect 23707 10016 24777 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 24765 10013 24777 10016
rect 24811 10013 24823 10047
rect 24765 10007 24823 10013
rect 27982 10004 27988 10056
rect 28040 10044 28046 10056
rect 28353 10047 28411 10053
rect 28353 10044 28365 10047
rect 28040 10016 28365 10044
rect 28040 10004 28046 10016
rect 28353 10013 28365 10016
rect 28399 10044 28411 10047
rect 28399 10016 28488 10044
rect 28399 10013 28411 10016
rect 28353 10007 28411 10013
rect 25130 9976 25136 9988
rect 20548 9948 22094 9976
rect 23032 9948 23612 9976
rect 23676 9948 25136 9976
rect 19429 9939 19487 9945
rect 20257 9911 20315 9917
rect 20257 9877 20269 9911
rect 20303 9908 20315 9911
rect 20898 9908 20904 9920
rect 20303 9880 20904 9908
rect 20303 9877 20315 9880
rect 20257 9871 20315 9877
rect 20898 9868 20904 9880
rect 20956 9868 20962 9920
rect 22066 9908 22094 9948
rect 22186 9908 22192 9920
rect 22066 9880 22192 9908
rect 22186 9868 22192 9880
rect 22244 9908 22250 9920
rect 23290 9908 23296 9920
rect 22244 9880 23296 9908
rect 22244 9868 22250 9880
rect 23290 9868 23296 9880
rect 23348 9868 23354 9920
rect 23474 9868 23480 9920
rect 23532 9908 23538 9920
rect 23676 9908 23704 9948
rect 25130 9936 25136 9948
rect 25188 9976 25194 9988
rect 26050 9976 26056 9988
rect 25188 9948 26056 9976
rect 25188 9936 25194 9948
rect 26050 9936 26056 9948
rect 26108 9936 26114 9988
rect 28460 9976 28488 10016
rect 28902 10004 28908 10056
rect 28960 10044 28966 10056
rect 29380 10044 29408 10084
rect 29546 10044 29552 10056
rect 28960 10016 29408 10044
rect 29507 10016 29552 10044
rect 28960 10004 28966 10016
rect 29546 10004 29552 10016
rect 29604 10004 29610 10056
rect 29733 9979 29791 9985
rect 29733 9976 29745 9979
rect 28460 9948 29745 9976
rect 29733 9945 29745 9948
rect 29779 9945 29791 9979
rect 29733 9939 29791 9945
rect 23842 9908 23848 9920
rect 23532 9880 23704 9908
rect 23803 9880 23848 9908
rect 23532 9868 23538 9880
rect 23842 9868 23848 9880
rect 23900 9868 23906 9920
rect 24578 9868 24584 9920
rect 24636 9908 24642 9920
rect 25774 9908 25780 9920
rect 24636 9880 25780 9908
rect 24636 9868 24642 9880
rect 25774 9868 25780 9880
rect 25832 9868 25838 9920
rect 26418 9908 26424 9920
rect 26379 9880 26424 9908
rect 26418 9868 26424 9880
rect 26476 9868 26482 9920
rect 28166 9868 28172 9920
rect 28224 9908 28230 9920
rect 28905 9911 28963 9917
rect 28905 9908 28917 9911
rect 28224 9880 28917 9908
rect 28224 9868 28230 9880
rect 28905 9877 28917 9880
rect 28951 9877 28963 9911
rect 29840 9908 29868 10084
rect 30561 10047 30619 10053
rect 30561 10013 30573 10047
rect 30607 10044 30619 10047
rect 30650 10044 30656 10056
rect 30607 10016 30656 10044
rect 30607 10013 30619 10016
rect 30561 10007 30619 10013
rect 30650 10004 30656 10016
rect 30708 10004 30714 10056
rect 30834 10053 30840 10056
rect 30828 10044 30840 10053
rect 30795 10016 30840 10044
rect 30828 10007 30840 10016
rect 30834 10004 30840 10007
rect 30892 10004 30898 10056
rect 42426 9976 42432 9988
rect 35866 9948 42432 9976
rect 35866 9908 35894 9948
rect 42426 9936 42432 9948
rect 42484 9976 42490 9988
rect 46842 9976 46848 9988
rect 42484 9948 46848 9976
rect 42484 9936 42490 9948
rect 46842 9936 46848 9948
rect 46900 9936 46906 9988
rect 29840 9880 35894 9908
rect 28905 9871 28963 9877
rect 1104 9818 48852 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 48852 9818
rect 1104 9744 48852 9766
rect 18046 9704 18052 9716
rect 17788 9676 18052 9704
rect 2958 9596 2964 9648
rect 3016 9636 3022 9648
rect 17788 9636 17816 9676
rect 18046 9664 18052 9676
rect 18104 9664 18110 9716
rect 20714 9664 20720 9716
rect 20772 9704 20778 9716
rect 20809 9707 20867 9713
rect 20809 9704 20821 9707
rect 20772 9676 20821 9704
rect 20772 9664 20778 9676
rect 20809 9673 20821 9676
rect 20855 9673 20867 9707
rect 20809 9667 20867 9673
rect 24394 9664 24400 9716
rect 24452 9704 24458 9716
rect 24489 9707 24547 9713
rect 24489 9704 24501 9707
rect 24452 9676 24501 9704
rect 24452 9664 24458 9676
rect 24489 9673 24501 9676
rect 24535 9673 24547 9707
rect 24489 9667 24547 9673
rect 28258 9664 28264 9716
rect 28316 9704 28322 9716
rect 29454 9704 29460 9716
rect 28316 9676 29460 9704
rect 28316 9664 28322 9676
rect 29454 9664 29460 9676
rect 29512 9664 29518 9716
rect 29641 9707 29699 9713
rect 29641 9673 29653 9707
rect 29687 9704 29699 9707
rect 29730 9704 29736 9716
rect 29687 9676 29736 9704
rect 29687 9673 29699 9676
rect 29641 9667 29699 9673
rect 29730 9664 29736 9676
rect 29788 9664 29794 9716
rect 21082 9636 21088 9648
rect 3016 9608 17816 9636
rect 17880 9608 21088 9636
rect 3016 9596 3022 9608
rect 17310 9528 17316 9580
rect 17368 9568 17374 9580
rect 17880 9577 17908 9608
rect 21082 9596 21088 9608
rect 21140 9596 21146 9648
rect 25958 9636 25964 9648
rect 23124 9608 25964 9636
rect 17865 9571 17923 9577
rect 17865 9568 17877 9571
rect 17368 9540 17877 9568
rect 17368 9528 17374 9540
rect 17865 9537 17877 9540
rect 17911 9537 17923 9571
rect 17865 9531 17923 9537
rect 18132 9571 18190 9577
rect 18132 9537 18144 9571
rect 18178 9568 18190 9571
rect 19058 9568 19064 9580
rect 18178 9540 19064 9568
rect 18178 9537 18190 9540
rect 18132 9531 18190 9537
rect 19058 9528 19064 9540
rect 19116 9528 19122 9580
rect 19242 9528 19248 9580
rect 19300 9568 19306 9580
rect 20441 9571 20499 9577
rect 20441 9568 20453 9571
rect 19300 9540 20453 9568
rect 19300 9528 19306 9540
rect 20441 9537 20453 9540
rect 20487 9537 20499 9571
rect 20441 9531 20499 9537
rect 20625 9571 20683 9577
rect 20625 9537 20637 9571
rect 20671 9568 20683 9571
rect 21910 9568 21916 9580
rect 20671 9540 21916 9568
rect 20671 9537 20683 9540
rect 20625 9531 20683 9537
rect 21910 9528 21916 9540
rect 21968 9528 21974 9580
rect 23124 9577 23152 9608
rect 25958 9596 25964 9608
rect 26016 9596 26022 9648
rect 26510 9636 26516 9648
rect 26160 9608 26516 9636
rect 23109 9571 23167 9577
rect 23109 9537 23121 9571
rect 23155 9537 23167 9571
rect 23109 9531 23167 9537
rect 23376 9571 23434 9577
rect 23376 9537 23388 9571
rect 23422 9568 23434 9571
rect 23842 9568 23848 9580
rect 23422 9540 23848 9568
rect 23422 9537 23434 9540
rect 23376 9531 23434 9537
rect 23842 9528 23848 9540
rect 23900 9528 23906 9580
rect 25685 9571 25743 9577
rect 25685 9570 25697 9571
rect 25608 9542 25697 9570
rect 25608 9432 25636 9542
rect 25685 9537 25697 9542
rect 25731 9537 25743 9571
rect 25685 9531 25743 9537
rect 25774 9528 25780 9580
rect 25832 9568 25838 9580
rect 25869 9571 25927 9577
rect 25869 9568 25881 9571
rect 25832 9540 25881 9568
rect 25832 9528 25838 9540
rect 25869 9537 25881 9540
rect 25915 9537 25927 9571
rect 26160 9568 26188 9608
rect 26510 9596 26516 9608
rect 26568 9596 26574 9648
rect 25869 9531 25927 9537
rect 25976 9540 26188 9568
rect 26237 9571 26295 9577
rect 25976 9509 26004 9540
rect 26237 9537 26249 9571
rect 26283 9568 26295 9571
rect 26418 9568 26424 9580
rect 26283 9540 26424 9568
rect 26283 9537 26295 9540
rect 26237 9531 26295 9537
rect 26418 9528 26424 9540
rect 26476 9528 26482 9580
rect 28353 9571 28411 9577
rect 28353 9537 28365 9571
rect 28399 9568 28411 9571
rect 28626 9568 28632 9580
rect 28399 9540 28632 9568
rect 28399 9537 28411 9540
rect 28353 9531 28411 9537
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29457 9571 29515 9577
rect 29457 9568 29469 9571
rect 29052 9540 29469 9568
rect 29052 9528 29058 9540
rect 29457 9537 29469 9540
rect 29503 9537 29515 9571
rect 29457 9531 29515 9537
rect 29641 9571 29699 9577
rect 29641 9537 29653 9571
rect 29687 9568 29699 9571
rect 29822 9568 29828 9580
rect 29687 9540 29828 9568
rect 29687 9537 29699 9540
rect 29641 9531 29699 9537
rect 29822 9528 29828 9540
rect 29880 9528 29886 9580
rect 25961 9503 26019 9509
rect 25961 9469 25973 9503
rect 26007 9469 26019 9503
rect 25961 9463 26019 9469
rect 26050 9460 26056 9512
rect 26108 9500 26114 9512
rect 28442 9500 28448 9512
rect 26108 9472 26153 9500
rect 28403 9472 28448 9500
rect 26108 9460 26114 9472
rect 28442 9460 28448 9472
rect 28500 9460 28506 9512
rect 28534 9460 28540 9512
rect 28592 9500 28598 9512
rect 28592 9472 28637 9500
rect 28592 9460 28598 9472
rect 26326 9432 26332 9444
rect 25608 9404 26332 9432
rect 26326 9392 26332 9404
rect 26384 9392 26390 9444
rect 27614 9392 27620 9444
rect 27672 9432 27678 9444
rect 27985 9435 28043 9441
rect 27985 9432 27997 9435
rect 27672 9404 27997 9432
rect 27672 9392 27678 9404
rect 27985 9401 27997 9404
rect 28031 9401 28043 9435
rect 27985 9395 28043 9401
rect 19245 9367 19303 9373
rect 19245 9333 19257 9367
rect 19291 9364 19303 9367
rect 19334 9364 19340 9376
rect 19291 9336 19340 9364
rect 19291 9333 19303 9336
rect 19245 9327 19303 9333
rect 19334 9324 19340 9336
rect 19392 9324 19398 9376
rect 26234 9324 26240 9376
rect 26292 9364 26298 9376
rect 26421 9367 26479 9373
rect 26421 9364 26433 9367
rect 26292 9336 26433 9364
rect 26292 9324 26298 9336
rect 26421 9333 26433 9336
rect 26467 9333 26479 9367
rect 26421 9327 26479 9333
rect 1104 9274 48852 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 48852 9274
rect 1104 9200 48852 9222
rect 20254 9160 20260 9172
rect 19904 9132 20260 9160
rect 17310 9024 17316 9036
rect 17271 8996 17316 9024
rect 17310 8984 17316 8996
rect 17368 8984 17374 9036
rect 19904 8965 19932 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 25774 9120 25780 9172
rect 25832 9160 25838 9172
rect 27338 9160 27344 9172
rect 25832 9132 27200 9160
rect 27299 9132 27344 9160
rect 25832 9120 25838 9132
rect 19978 9052 19984 9104
rect 20036 9052 20042 9104
rect 19996 9024 20024 9052
rect 25958 9024 25964 9036
rect 19996 8996 20208 9024
rect 25919 8996 25964 9024
rect 20180 8968 20208 8996
rect 25958 8984 25964 8996
rect 26016 8984 26022 9036
rect 27172 9024 27200 9132
rect 27338 9120 27344 9132
rect 27396 9120 27402 9172
rect 27430 9120 27436 9172
rect 27488 9160 27494 9172
rect 32582 9160 32588 9172
rect 27488 9132 32588 9160
rect 27488 9120 27494 9132
rect 32582 9120 32588 9132
rect 32640 9120 32646 9172
rect 28534 9052 28540 9104
rect 28592 9092 28598 9104
rect 30098 9092 30104 9104
rect 28592 9064 30104 9092
rect 28592 9052 28598 9064
rect 30098 9052 30104 9064
rect 30156 9052 30162 9104
rect 28258 9024 28264 9036
rect 27172 8996 28264 9024
rect 28258 8984 28264 8996
rect 28316 9024 28322 9036
rect 28316 8996 28396 9024
rect 28316 8984 28322 8996
rect 19797 8959 19855 8965
rect 19797 8925 19809 8959
rect 19843 8925 19855 8959
rect 19797 8919 19855 8925
rect 19889 8959 19947 8965
rect 19889 8925 19901 8959
rect 19935 8925 19947 8959
rect 19889 8919 19947 8925
rect 17580 8891 17638 8897
rect 17580 8857 17592 8891
rect 17626 8888 17638 8891
rect 19521 8891 19579 8897
rect 19521 8888 19533 8891
rect 17626 8860 19533 8888
rect 17626 8857 17638 8860
rect 17580 8851 17638 8857
rect 19521 8857 19533 8860
rect 19567 8857 19579 8891
rect 19812 8888 19840 8919
rect 19978 8916 19984 8968
rect 20036 8956 20042 8968
rect 20036 8928 20081 8956
rect 20036 8916 20042 8928
rect 20162 8916 20168 8968
rect 20220 8956 20226 8968
rect 20625 8959 20683 8965
rect 20220 8928 20313 8956
rect 20220 8916 20226 8928
rect 20625 8925 20637 8959
rect 20671 8956 20683 8959
rect 20714 8956 20720 8968
rect 20671 8928 20720 8956
rect 20671 8925 20683 8928
rect 20625 8919 20683 8925
rect 20714 8916 20720 8928
rect 20772 8916 20778 8968
rect 20898 8965 20904 8968
rect 20892 8956 20904 8965
rect 20859 8928 20904 8956
rect 20892 8919 20904 8928
rect 20898 8916 20904 8919
rect 20956 8916 20962 8968
rect 26234 8965 26240 8968
rect 26228 8956 26240 8965
rect 26195 8928 26240 8956
rect 26228 8919 26240 8928
rect 26234 8916 26240 8919
rect 26292 8916 26298 8968
rect 28166 8956 28172 8968
rect 28127 8928 28172 8956
rect 28166 8916 28172 8928
rect 28224 8916 28230 8968
rect 28368 8965 28396 8996
rect 28442 8984 28448 9036
rect 28500 9024 28506 9036
rect 29270 9024 29276 9036
rect 28500 8996 29276 9024
rect 28500 8984 28506 8996
rect 29270 8984 29276 8996
rect 29328 9024 29334 9036
rect 29730 9024 29736 9036
rect 29328 8996 29736 9024
rect 29328 8984 29334 8996
rect 29730 8984 29736 8996
rect 29788 8984 29794 9036
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8925 28411 8959
rect 28534 8956 28540 8968
rect 28495 8928 28540 8956
rect 28353 8919 28411 8925
rect 28534 8916 28540 8928
rect 28592 8916 28598 8968
rect 28626 8916 28632 8968
rect 28684 8956 28690 8968
rect 28721 8959 28779 8965
rect 28721 8956 28733 8959
rect 28684 8928 28733 8956
rect 28684 8916 28690 8928
rect 28721 8925 28733 8928
rect 28767 8925 28779 8959
rect 28721 8919 28779 8925
rect 20806 8888 20812 8900
rect 19812 8860 20812 8888
rect 19521 8851 19579 8857
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 26878 8848 26884 8900
rect 26936 8888 26942 8900
rect 28644 8888 28672 8916
rect 26936 8860 28672 8888
rect 26936 8848 26942 8860
rect 28810 8848 28816 8900
rect 28868 8888 28874 8900
rect 30742 8888 30748 8900
rect 28868 8860 30748 8888
rect 28868 8848 28874 8860
rect 30742 8848 30748 8860
rect 30800 8848 30806 8900
rect 47946 8888 47952 8900
rect 47907 8860 47952 8888
rect 47946 8848 47952 8860
rect 48004 8848 48010 8900
rect 18693 8823 18751 8829
rect 18693 8789 18705 8823
rect 18739 8820 18751 8823
rect 18874 8820 18880 8832
rect 18739 8792 18880 8820
rect 18739 8789 18751 8792
rect 18693 8783 18751 8789
rect 18874 8780 18880 8792
rect 18932 8780 18938 8832
rect 20714 8780 20720 8832
rect 20772 8820 20778 8832
rect 21082 8820 21088 8832
rect 20772 8792 21088 8820
rect 20772 8780 20778 8792
rect 21082 8780 21088 8792
rect 21140 8780 21146 8832
rect 21910 8780 21916 8832
rect 21968 8820 21974 8832
rect 22005 8823 22063 8829
rect 22005 8820 22017 8823
rect 21968 8792 22017 8820
rect 21968 8780 21974 8792
rect 22005 8789 22017 8792
rect 22051 8789 22063 8823
rect 28902 8820 28908 8832
rect 28863 8792 28908 8820
rect 22005 8783 22063 8789
rect 28902 8780 28908 8792
rect 28960 8780 28966 8832
rect 38286 8780 38292 8832
rect 38344 8820 38350 8832
rect 48041 8823 48099 8829
rect 48041 8820 48053 8823
rect 38344 8792 48053 8820
rect 38344 8780 38350 8792
rect 48041 8789 48053 8792
rect 48087 8789 48099 8823
rect 48041 8783 48099 8789
rect 1104 8730 48852 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 48852 8730
rect 1104 8656 48852 8678
rect 27522 8576 27528 8628
rect 27580 8616 27586 8628
rect 29730 8616 29736 8628
rect 27580 8588 29040 8616
rect 29691 8588 29736 8616
rect 27580 8576 27586 8588
rect 19334 8548 19340 8560
rect 18524 8520 19340 8548
rect 1854 8480 1860 8492
rect 1815 8452 1860 8480
rect 1854 8440 1860 8452
rect 1912 8440 1918 8492
rect 18524 8489 18552 8520
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 28353 8483 28411 8489
rect 28353 8449 28365 8483
rect 28399 8449 28411 8483
rect 28353 8443 28411 8449
rect 28620 8483 28678 8489
rect 28620 8449 28632 8483
rect 28666 8480 28678 8483
rect 28902 8480 28908 8492
rect 28666 8452 28908 8480
rect 28666 8449 28678 8452
rect 28620 8443 28678 8449
rect 18690 8412 18696 8424
rect 18651 8384 18696 8412
rect 18690 8372 18696 8384
rect 18748 8372 18754 8424
rect 19426 8412 19432 8424
rect 19387 8384 19432 8412
rect 19426 8372 19432 8384
rect 19484 8372 19490 8424
rect 20806 8372 20812 8424
rect 20864 8412 20870 8424
rect 21818 8412 21824 8424
rect 20864 8384 21824 8412
rect 20864 8372 20870 8384
rect 21818 8372 21824 8384
rect 21876 8412 21882 8424
rect 26418 8412 26424 8424
rect 21876 8384 26424 8412
rect 21876 8372 21882 8384
rect 26418 8372 26424 8384
rect 26476 8372 26482 8424
rect 2133 8347 2191 8353
rect 2133 8313 2145 8347
rect 2179 8344 2191 8347
rect 16666 8344 16672 8356
rect 2179 8316 16672 8344
rect 2179 8313 2191 8316
rect 2133 8307 2191 8313
rect 16666 8304 16672 8316
rect 16724 8304 16730 8356
rect 20162 8304 20168 8356
rect 20220 8344 20226 8356
rect 27430 8344 27436 8356
rect 20220 8316 27436 8344
rect 20220 8304 20226 8316
rect 27430 8304 27436 8316
rect 27488 8304 27494 8356
rect 28368 8276 28396 8443
rect 28902 8440 28908 8452
rect 28960 8440 28966 8492
rect 29012 8480 29040 8588
rect 29730 8576 29736 8588
rect 29788 8576 29794 8628
rect 30742 8576 30748 8628
rect 30800 8616 30806 8628
rect 47857 8619 47915 8625
rect 47857 8616 47869 8619
rect 30800 8588 47869 8616
rect 30800 8576 30806 8588
rect 47857 8585 47869 8588
rect 47903 8585 47915 8619
rect 47857 8579 47915 8585
rect 30466 8480 30472 8492
rect 29012 8452 30328 8480
rect 30427 8452 30472 8480
rect 30300 8412 30328 8452
rect 30466 8440 30472 8452
rect 30524 8440 30530 8492
rect 30561 8483 30619 8489
rect 30561 8449 30573 8483
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 30653 8483 30711 8489
rect 30653 8449 30665 8483
rect 30699 8449 30711 8483
rect 30653 8443 30711 8449
rect 30837 8483 30895 8489
rect 30837 8449 30849 8483
rect 30883 8480 30895 8483
rect 32582 8480 32588 8492
rect 30883 8452 32588 8480
rect 30883 8449 30895 8452
rect 30837 8443 30895 8449
rect 30576 8412 30604 8443
rect 30300 8384 30604 8412
rect 30668 8412 30696 8443
rect 32582 8440 32588 8452
rect 32640 8440 32646 8492
rect 47762 8480 47768 8492
rect 47723 8452 47768 8480
rect 47762 8440 47768 8452
rect 47820 8440 47826 8492
rect 31846 8412 31852 8424
rect 30668 8384 31852 8412
rect 31846 8372 31852 8384
rect 31904 8372 31910 8424
rect 30650 8344 30656 8356
rect 29288 8316 30656 8344
rect 29288 8276 29316 8316
rect 30650 8304 30656 8316
rect 30708 8304 30714 8356
rect 30190 8276 30196 8288
rect 28368 8248 29316 8276
rect 30151 8248 30196 8276
rect 30190 8236 30196 8248
rect 30248 8236 30254 8288
rect 1104 8186 48852 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 48852 8186
rect 1104 8112 48852 8134
rect 18601 8075 18659 8081
rect 18601 8041 18613 8075
rect 18647 8072 18659 8075
rect 18690 8072 18696 8084
rect 18647 8044 18696 8072
rect 18647 8041 18659 8044
rect 18601 8035 18659 8041
rect 18690 8032 18696 8044
rect 18748 8032 18754 8084
rect 19797 8075 19855 8081
rect 19797 8041 19809 8075
rect 19843 8072 19855 8075
rect 19978 8072 19984 8084
rect 19843 8044 19984 8072
rect 19843 8041 19855 8044
rect 19797 8035 19855 8041
rect 19978 8032 19984 8044
rect 20036 8032 20042 8084
rect 20714 8032 20720 8084
rect 20772 8072 20778 8084
rect 21726 8072 21732 8084
rect 20772 8044 21732 8072
rect 20772 8032 20778 8044
rect 21726 8032 21732 8044
rect 21784 8072 21790 8084
rect 23842 8072 23848 8084
rect 21784 8044 23848 8072
rect 21784 8032 21790 8044
rect 23842 8032 23848 8044
rect 23900 8032 23906 8084
rect 31846 8072 31852 8084
rect 29564 8044 30788 8072
rect 31807 8044 31852 8072
rect 21358 7964 21364 8016
rect 21416 7964 21422 8016
rect 22094 8004 22100 8016
rect 22020 7976 22100 8004
rect 16482 7896 16488 7948
rect 16540 7936 16546 7948
rect 21376 7936 21404 7964
rect 16540 7908 21220 7936
rect 16540 7896 16546 7908
rect 18509 7871 18567 7877
rect 18509 7837 18521 7871
rect 18555 7837 18567 7871
rect 18509 7831 18567 7837
rect 1854 7800 1860 7812
rect 1815 7772 1860 7800
rect 1854 7760 1860 7772
rect 1912 7760 1918 7812
rect 18524 7800 18552 7831
rect 18874 7828 18880 7880
rect 18932 7868 18938 7880
rect 21192 7877 21220 7908
rect 21284 7908 21404 7936
rect 21284 7877 21312 7908
rect 19613 7871 19671 7877
rect 19613 7868 19625 7871
rect 18932 7840 19625 7868
rect 18932 7828 18938 7840
rect 19613 7837 19625 7840
rect 19659 7837 19671 7871
rect 19613 7831 19671 7837
rect 21177 7871 21235 7877
rect 21177 7837 21189 7871
rect 21223 7837 21235 7871
rect 21177 7831 21235 7837
rect 21266 7871 21324 7877
rect 21266 7837 21278 7871
rect 21312 7837 21324 7871
rect 21266 7831 21324 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21545 7871 21603 7877
rect 21545 7837 21557 7871
rect 21591 7868 21603 7871
rect 21726 7868 21732 7880
rect 21591 7840 21732 7868
rect 21591 7837 21603 7840
rect 21545 7831 21603 7837
rect 19242 7800 19248 7812
rect 18524 7772 19248 7800
rect 19242 7760 19248 7772
rect 19300 7760 19306 7812
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 19392 7772 19441 7800
rect 19392 7760 19398 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 21376 7800 21404 7831
rect 21726 7828 21732 7840
rect 21784 7828 21790 7880
rect 22020 7877 22048 7976
rect 22094 7964 22100 7976
rect 22152 8004 22158 8016
rect 22278 8004 22284 8016
rect 22152 7976 22284 8004
rect 22152 7964 22158 7976
rect 22278 7964 22284 7976
rect 22336 7964 22342 8016
rect 23658 8004 23664 8016
rect 23584 7976 23664 8004
rect 22005 7871 22063 7877
rect 22005 7837 22017 7871
rect 22051 7837 22063 7871
rect 22005 7831 22063 7837
rect 22186 7828 22192 7880
rect 22244 7868 22250 7880
rect 22244 7840 22289 7868
rect 22244 7828 22250 7840
rect 22646 7828 22652 7880
rect 22704 7868 22710 7880
rect 23584 7877 23612 7976
rect 23658 7964 23664 7976
rect 23716 7964 23722 8016
rect 24765 7939 24823 7945
rect 24765 7936 24777 7939
rect 23676 7908 24777 7936
rect 23676 7877 23704 7908
rect 24765 7905 24777 7908
rect 24811 7905 24823 7939
rect 28077 7939 28135 7945
rect 28077 7936 28089 7939
rect 24765 7899 24823 7905
rect 27080 7908 28089 7936
rect 23477 7871 23535 7877
rect 23477 7868 23489 7871
rect 22704 7840 23489 7868
rect 22704 7828 22710 7840
rect 23477 7837 23489 7840
rect 23523 7837 23535 7871
rect 23477 7831 23535 7837
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 23661 7871 23719 7877
rect 23661 7837 23673 7871
rect 23707 7837 23719 7871
rect 23842 7868 23848 7880
rect 23803 7840 23848 7868
rect 23661 7831 23719 7837
rect 23842 7828 23848 7840
rect 23900 7828 23906 7880
rect 24581 7871 24639 7877
rect 24581 7837 24593 7871
rect 24627 7868 24639 7871
rect 26878 7868 26884 7880
rect 24627 7840 26884 7868
rect 24627 7837 24639 7840
rect 24581 7831 24639 7837
rect 26878 7828 26884 7840
rect 26936 7828 26942 7880
rect 27080 7877 27108 7908
rect 28077 7905 28089 7908
rect 28123 7905 28135 7939
rect 28077 7899 28135 7905
rect 26973 7871 27031 7877
rect 26973 7837 26985 7871
rect 27019 7837 27031 7871
rect 26973 7831 27031 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27249 7871 27307 7877
rect 27249 7837 27261 7871
rect 27295 7868 27307 7871
rect 27430 7868 27436 7880
rect 27295 7840 27436 7868
rect 27295 7837 27307 7840
rect 27249 7831 27307 7837
rect 22094 7800 22100 7812
rect 21376 7772 22100 7800
rect 19429 7763 19487 7769
rect 22094 7760 22100 7772
rect 22152 7760 22158 7812
rect 22278 7760 22284 7812
rect 22336 7800 22342 7812
rect 24397 7803 24455 7809
rect 24397 7800 24409 7803
rect 22336 7772 24409 7800
rect 22336 7760 22342 7772
rect 24397 7769 24409 7772
rect 24443 7769 24455 7803
rect 26988 7800 27016 7831
rect 27430 7828 27436 7840
rect 27488 7828 27494 7880
rect 29564 7868 29592 8044
rect 27724 7840 29592 7868
rect 29641 7871 29699 7877
rect 27522 7800 27528 7812
rect 26988 7772 27528 7800
rect 24397 7763 24455 7769
rect 27522 7760 27528 7772
rect 27580 7760 27586 7812
rect 27724 7809 27752 7840
rect 29641 7837 29653 7871
rect 29687 7868 29699 7871
rect 30650 7868 30656 7880
rect 29687 7840 30656 7868
rect 29687 7837 29699 7840
rect 29641 7831 29699 7837
rect 30650 7828 30656 7840
rect 30708 7828 30714 7880
rect 30760 7868 30788 8044
rect 31846 8032 31852 8044
rect 31904 8032 31910 8084
rect 31481 7871 31539 7877
rect 31481 7868 31493 7871
rect 30760 7840 31493 7868
rect 31481 7837 31493 7840
rect 31527 7837 31539 7871
rect 31481 7831 31539 7837
rect 27709 7803 27767 7809
rect 27709 7769 27721 7803
rect 27755 7769 27767 7803
rect 27709 7763 27767 7769
rect 27893 7803 27951 7809
rect 27893 7769 27905 7803
rect 27939 7800 27951 7803
rect 28258 7800 28264 7812
rect 27939 7772 28264 7800
rect 27939 7769 27951 7772
rect 27893 7763 27951 7769
rect 2133 7735 2191 7741
rect 2133 7701 2145 7735
rect 2179 7732 2191 7735
rect 18966 7732 18972 7744
rect 2179 7704 18972 7732
rect 2179 7701 2191 7704
rect 2133 7695 2191 7701
rect 18966 7692 18972 7704
rect 19024 7692 19030 7744
rect 20898 7732 20904 7744
rect 20859 7704 20904 7732
rect 20898 7692 20904 7704
rect 20956 7692 20962 7744
rect 21450 7692 21456 7744
rect 21508 7732 21514 7744
rect 22373 7735 22431 7741
rect 22373 7732 22385 7735
rect 21508 7704 22385 7732
rect 21508 7692 21514 7704
rect 22373 7701 22385 7704
rect 22419 7701 22431 7735
rect 22373 7695 22431 7701
rect 23201 7735 23259 7741
rect 23201 7701 23213 7735
rect 23247 7732 23259 7735
rect 24486 7732 24492 7744
rect 23247 7704 24492 7732
rect 23247 7701 23259 7704
rect 23201 7695 23259 7701
rect 24486 7692 24492 7704
rect 24544 7692 24550 7744
rect 26602 7732 26608 7744
rect 26563 7704 26608 7732
rect 26602 7692 26608 7704
rect 26660 7692 26666 7744
rect 26970 7692 26976 7744
rect 27028 7732 27034 7744
rect 27724 7732 27752 7763
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 29908 7803 29966 7809
rect 29908 7769 29920 7803
rect 29954 7800 29966 7803
rect 30190 7800 30196 7812
rect 29954 7772 30196 7800
rect 29954 7769 29966 7772
rect 29908 7763 29966 7769
rect 30190 7760 30196 7772
rect 30248 7760 30254 7812
rect 31665 7803 31723 7809
rect 31665 7769 31677 7803
rect 31711 7769 31723 7803
rect 31665 7763 31723 7769
rect 27028 7704 27752 7732
rect 27028 7692 27034 7704
rect 29638 7692 29644 7744
rect 29696 7732 29702 7744
rect 31021 7735 31079 7741
rect 31021 7732 31033 7735
rect 29696 7704 31033 7732
rect 29696 7692 29702 7704
rect 31021 7701 31033 7704
rect 31067 7732 31079 7735
rect 31680 7732 31708 7763
rect 31067 7704 31708 7732
rect 31067 7701 31079 7704
rect 31021 7695 31079 7701
rect 1104 7642 48852 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 48852 7642
rect 1104 7568 48852 7590
rect 22186 7488 22192 7540
rect 22244 7528 22250 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 22244 7500 23213 7528
rect 22244 7488 22250 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 23201 7491 23259 7497
rect 25222 7488 25228 7540
rect 25280 7528 25286 7540
rect 25280 7500 41414 7528
rect 25280 7488 25286 7500
rect 19242 7420 19248 7472
rect 19300 7460 19306 7472
rect 19300 7432 26280 7460
rect 19300 7420 19306 7432
rect 18874 7392 18880 7404
rect 18835 7364 18880 7392
rect 18874 7352 18880 7364
rect 18932 7352 18938 7404
rect 20806 7352 20812 7404
rect 20864 7392 20870 7404
rect 22077 7395 22135 7401
rect 22077 7392 22089 7395
rect 20864 7364 22089 7392
rect 20864 7352 20870 7364
rect 22077 7361 22089 7364
rect 22123 7361 22135 7395
rect 22077 7355 22135 7361
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 26252 7401 26280 7432
rect 26602 7420 26608 7472
rect 26660 7460 26666 7472
rect 27218 7463 27276 7469
rect 27218 7460 27230 7463
rect 26660 7432 27230 7460
rect 26660 7420 26666 7432
rect 27218 7429 27230 7432
rect 27264 7429 27276 7463
rect 27218 7423 27276 7429
rect 23917 7395 23975 7401
rect 23917 7392 23929 7395
rect 23808 7364 23929 7392
rect 23808 7352 23814 7364
rect 23917 7361 23929 7364
rect 23963 7361 23975 7395
rect 23917 7355 23975 7361
rect 26237 7395 26295 7401
rect 26237 7361 26249 7395
rect 26283 7392 26295 7395
rect 27798 7392 27804 7404
rect 26283 7364 27804 7392
rect 26283 7361 26295 7364
rect 26237 7355 26295 7361
rect 27798 7352 27804 7364
rect 27856 7352 27862 7404
rect 29638 7392 29644 7404
rect 29599 7364 29644 7392
rect 29638 7352 29644 7364
rect 29696 7352 29702 7404
rect 41386 7392 41414 7500
rect 45738 7392 45744 7404
rect 41386 7364 45744 7392
rect 45738 7352 45744 7364
rect 45796 7392 45802 7404
rect 46661 7395 46719 7401
rect 46661 7392 46673 7395
rect 45796 7364 46673 7392
rect 45796 7352 45802 7364
rect 46661 7361 46673 7364
rect 46707 7361 46719 7395
rect 46661 7355 46719 7361
rect 19061 7327 19119 7333
rect 19061 7293 19073 7327
rect 19107 7324 19119 7327
rect 19334 7324 19340 7336
rect 19107 7296 19340 7324
rect 19107 7293 19119 7296
rect 19061 7287 19119 7293
rect 19334 7284 19340 7296
rect 19392 7284 19398 7336
rect 19429 7327 19487 7333
rect 19429 7293 19441 7327
rect 19475 7293 19487 7327
rect 19429 7287 19487 7293
rect 18690 7216 18696 7268
rect 18748 7256 18754 7268
rect 19444 7256 19472 7287
rect 21082 7284 21088 7336
rect 21140 7324 21146 7336
rect 21821 7327 21879 7333
rect 21821 7324 21833 7327
rect 21140 7296 21833 7324
rect 21140 7284 21146 7296
rect 21821 7293 21833 7296
rect 21867 7293 21879 7327
rect 21821 7287 21879 7293
rect 23661 7327 23719 7333
rect 23661 7293 23673 7327
rect 23707 7293 23719 7327
rect 23661 7287 23719 7293
rect 18748 7228 19472 7256
rect 18748 7216 18754 7228
rect 2038 7188 2044 7200
rect 1999 7160 2044 7188
rect 2038 7148 2044 7160
rect 2096 7148 2102 7200
rect 23676 7188 23704 7287
rect 25958 7284 25964 7336
rect 26016 7324 26022 7336
rect 26973 7327 27031 7333
rect 26973 7324 26985 7327
rect 26016 7296 26985 7324
rect 26016 7284 26022 7296
rect 26973 7293 26985 7296
rect 27019 7293 27031 7327
rect 29822 7324 29828 7336
rect 29783 7296 29828 7324
rect 26973 7287 27031 7293
rect 29822 7284 29828 7296
rect 29880 7284 29886 7336
rect 30101 7327 30159 7333
rect 30101 7293 30113 7327
rect 30147 7293 30159 7327
rect 30101 7287 30159 7293
rect 29638 7216 29644 7268
rect 29696 7256 29702 7268
rect 30116 7256 30144 7287
rect 29696 7228 30144 7256
rect 29696 7216 29702 7228
rect 24946 7188 24952 7200
rect 23676 7160 24952 7188
rect 24946 7148 24952 7160
rect 25004 7148 25010 7200
rect 25038 7148 25044 7200
rect 25096 7188 25102 7200
rect 26329 7191 26387 7197
rect 25096 7160 25141 7188
rect 25096 7148 25102 7160
rect 26329 7157 26341 7191
rect 26375 7188 26387 7191
rect 26694 7188 26700 7200
rect 26375 7160 26700 7188
rect 26375 7157 26387 7160
rect 26329 7151 26387 7157
rect 26694 7148 26700 7160
rect 26752 7148 26758 7200
rect 28258 7148 28264 7200
rect 28316 7188 28322 7200
rect 28353 7191 28411 7197
rect 28353 7188 28365 7191
rect 28316 7160 28365 7188
rect 28316 7148 28322 7160
rect 28353 7157 28365 7160
rect 28399 7157 28411 7191
rect 28353 7151 28411 7157
rect 46474 7148 46480 7200
rect 46532 7188 46538 7200
rect 46753 7191 46811 7197
rect 46753 7188 46765 7191
rect 46532 7160 46765 7188
rect 46532 7148 46538 7160
rect 46753 7157 46765 7160
rect 46799 7157 46811 7191
rect 47762 7188 47768 7200
rect 47723 7160 47768 7188
rect 46753 7151 46811 7157
rect 47762 7148 47768 7160
rect 47820 7148 47826 7200
rect 1104 7098 48852 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 48852 7098
rect 1104 7024 48852 7046
rect 21818 6944 21824 6996
rect 21876 6984 21882 6996
rect 22094 6984 22100 6996
rect 21876 6956 22100 6984
rect 21876 6944 21882 6956
rect 22094 6944 22100 6956
rect 22152 6984 22158 6996
rect 22465 6987 22523 6993
rect 22465 6984 22477 6987
rect 22152 6956 22477 6984
rect 22152 6944 22158 6956
rect 22465 6953 22477 6956
rect 22511 6953 22523 6987
rect 22465 6947 22523 6953
rect 25777 6987 25835 6993
rect 25777 6953 25789 6987
rect 25823 6984 25835 6987
rect 26878 6984 26884 6996
rect 25823 6956 26884 6984
rect 25823 6953 25835 6956
rect 25777 6947 25835 6953
rect 26878 6944 26884 6956
rect 26936 6944 26942 6996
rect 29822 6984 29828 6996
rect 29783 6956 29828 6984
rect 29822 6944 29828 6956
rect 29880 6944 29886 6996
rect 1397 6851 1455 6857
rect 1397 6817 1409 6851
rect 1443 6848 1455 6851
rect 2038 6848 2044 6860
rect 1443 6820 2044 6848
rect 1443 6817 1455 6820
rect 1397 6811 1455 6817
rect 2038 6808 2044 6820
rect 2096 6808 2102 6860
rect 2774 6848 2780 6860
rect 2735 6820 2780 6848
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 19334 6848 19340 6860
rect 19295 6820 19340 6848
rect 19334 6808 19340 6820
rect 19392 6808 19398 6860
rect 19981 6851 20039 6857
rect 19981 6817 19993 6851
rect 20027 6848 20039 6851
rect 20806 6848 20812 6860
rect 20027 6820 20812 6848
rect 20027 6817 20039 6820
rect 19981 6811 20039 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 21082 6848 21088 6860
rect 21043 6820 21088 6848
rect 21082 6808 21088 6820
rect 21140 6808 21146 6860
rect 23201 6851 23259 6857
rect 23201 6817 23213 6851
rect 23247 6848 23259 6851
rect 23750 6848 23756 6860
rect 23247 6820 23756 6848
rect 23247 6817 23259 6820
rect 23201 6811 23259 6817
rect 23750 6808 23756 6820
rect 23808 6808 23814 6860
rect 26694 6848 26700 6860
rect 26655 6820 26700 6848
rect 26694 6808 26700 6820
rect 26752 6808 26758 6860
rect 26970 6848 26976 6860
rect 26931 6820 26976 6848
rect 26970 6808 26976 6820
rect 27028 6808 27034 6860
rect 37090 6808 37096 6860
rect 37148 6848 37154 6860
rect 45646 6848 45652 6860
rect 37148 6820 45652 6848
rect 37148 6808 37154 6820
rect 45646 6808 45652 6820
rect 45704 6808 45710 6860
rect 46474 6848 46480 6860
rect 46435 6820 46480 6848
rect 46474 6808 46480 6820
rect 46532 6808 46538 6860
rect 48130 6848 48136 6860
rect 48091 6820 48136 6848
rect 48130 6808 48136 6820
rect 48188 6808 48194 6860
rect 19242 6780 19248 6792
rect 19203 6752 19248 6780
rect 19242 6740 19248 6752
rect 19300 6740 19306 6792
rect 20257 6783 20315 6789
rect 20257 6749 20269 6783
rect 20303 6749 20315 6783
rect 20257 6743 20315 6749
rect 20349 6783 20407 6789
rect 20349 6749 20361 6783
rect 20395 6749 20407 6783
rect 20349 6743 20407 6749
rect 20441 6783 20499 6789
rect 20441 6749 20453 6783
rect 20487 6749 20499 6783
rect 20441 6743 20499 6749
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6780 20683 6783
rect 20714 6780 20720 6792
rect 20671 6752 20720 6780
rect 20671 6749 20683 6752
rect 20625 6743 20683 6749
rect 1581 6715 1639 6721
rect 1581 6681 1593 6715
rect 1627 6712 1639 6715
rect 2222 6712 2228 6724
rect 1627 6684 2228 6712
rect 1627 6681 1639 6684
rect 1581 6675 1639 6681
rect 2222 6672 2228 6684
rect 2280 6672 2286 6724
rect 15194 6672 15200 6724
rect 15252 6712 15258 6724
rect 20272 6712 20300 6743
rect 15252 6684 20300 6712
rect 15252 6672 15258 6684
rect 20364 6644 20392 6743
rect 20456 6712 20484 6743
rect 20714 6740 20720 6752
rect 20772 6740 20778 6792
rect 20898 6740 20904 6792
rect 20956 6780 20962 6792
rect 21341 6783 21399 6789
rect 21341 6780 21353 6783
rect 20956 6752 21353 6780
rect 20956 6740 20962 6752
rect 21341 6749 21353 6752
rect 21387 6749 21399 6783
rect 21341 6743 21399 6749
rect 23382 6740 23388 6792
rect 23440 6789 23446 6792
rect 23440 6783 23489 6789
rect 23440 6749 23443 6783
rect 23477 6749 23489 6783
rect 23566 6780 23572 6792
rect 23527 6752 23572 6780
rect 23440 6743 23489 6749
rect 23440 6740 23446 6743
rect 23566 6740 23572 6752
rect 23624 6740 23630 6792
rect 23658 6740 23664 6792
rect 23716 6780 23722 6792
rect 23845 6783 23903 6789
rect 23716 6752 23761 6780
rect 23716 6740 23722 6752
rect 23845 6749 23857 6783
rect 23891 6780 23903 6783
rect 24026 6780 24032 6792
rect 23891 6752 24032 6780
rect 23891 6749 23903 6752
rect 23845 6743 23903 6749
rect 24026 6740 24032 6752
rect 24084 6740 24090 6792
rect 24397 6783 24455 6789
rect 24397 6749 24409 6783
rect 24443 6780 24455 6783
rect 24946 6780 24952 6792
rect 24443 6752 24952 6780
rect 24443 6749 24455 6752
rect 24397 6743 24455 6749
rect 24946 6740 24952 6752
rect 25004 6780 25010 6792
rect 25958 6780 25964 6792
rect 25004 6752 25964 6780
rect 25004 6740 25010 6752
rect 25958 6740 25964 6752
rect 26016 6740 26022 6792
rect 26513 6783 26571 6789
rect 26513 6749 26525 6783
rect 26559 6749 26571 6783
rect 26513 6743 26571 6749
rect 21450 6712 21456 6724
rect 20456 6684 21456 6712
rect 21450 6672 21456 6684
rect 21508 6672 21514 6724
rect 24486 6672 24492 6724
rect 24544 6712 24550 6724
rect 24642 6715 24700 6721
rect 24642 6712 24654 6715
rect 24544 6684 24654 6712
rect 24544 6672 24550 6684
rect 24642 6681 24654 6684
rect 24688 6681 24700 6715
rect 26528 6712 26556 6743
rect 27890 6740 27896 6792
rect 27948 6780 27954 6792
rect 29733 6783 29791 6789
rect 29733 6780 29745 6783
rect 27948 6752 29745 6780
rect 27948 6740 27954 6752
rect 29733 6749 29745 6752
rect 29779 6749 29791 6783
rect 29733 6743 29791 6749
rect 46293 6783 46351 6789
rect 46293 6749 46305 6783
rect 46339 6749 46351 6783
rect 46293 6743 46351 6749
rect 28258 6712 28264 6724
rect 26528 6684 28264 6712
rect 24642 6675 24700 6681
rect 28258 6672 28264 6684
rect 28316 6672 28322 6724
rect 37182 6672 37188 6724
rect 37240 6712 37246 6724
rect 45554 6712 45560 6724
rect 37240 6684 45560 6712
rect 37240 6672 37246 6684
rect 45554 6672 45560 6684
rect 45612 6672 45618 6724
rect 46308 6712 46336 6743
rect 47762 6712 47768 6724
rect 46308 6684 47768 6712
rect 47762 6672 47768 6684
rect 47820 6672 47826 6724
rect 21542 6644 21548 6656
rect 20364 6616 21548 6644
rect 21542 6604 21548 6616
rect 21600 6644 21606 6656
rect 23566 6644 23572 6656
rect 21600 6616 23572 6644
rect 21600 6604 21606 6616
rect 23566 6604 23572 6616
rect 23624 6604 23630 6656
rect 1104 6554 48852 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 48852 6554
rect 1104 6480 48852 6502
rect 2222 6440 2228 6452
rect 2183 6412 2228 6440
rect 2222 6400 2228 6412
rect 2280 6400 2286 6452
rect 22186 6440 22192 6452
rect 22147 6412 22192 6440
rect 22186 6400 22192 6412
rect 22244 6400 22250 6452
rect 23477 6443 23535 6449
rect 23477 6409 23489 6443
rect 23523 6440 23535 6443
rect 23658 6440 23664 6452
rect 23523 6412 23664 6440
rect 23523 6409 23535 6412
rect 23477 6403 23535 6409
rect 23658 6400 23664 6412
rect 23716 6400 23722 6452
rect 38654 6440 38660 6452
rect 26206 6412 38660 6440
rect 22005 6375 22063 6381
rect 22005 6341 22017 6375
rect 22051 6372 22063 6375
rect 22094 6372 22100 6384
rect 22051 6344 22100 6372
rect 22051 6341 22063 6344
rect 22005 6335 22063 6341
rect 22094 6332 22100 6344
rect 22152 6332 22158 6384
rect 23293 6375 23351 6381
rect 23293 6341 23305 6375
rect 23339 6372 23351 6375
rect 25038 6372 25044 6384
rect 23339 6344 25044 6372
rect 23339 6341 23351 6344
rect 23293 6335 23351 6341
rect 25038 6332 25044 6344
rect 25096 6332 25102 6384
rect 2130 6304 2136 6316
rect 2091 6276 2136 6304
rect 2130 6264 2136 6276
rect 2188 6264 2194 6316
rect 21821 6307 21879 6313
rect 21821 6273 21833 6307
rect 21867 6273 21879 6307
rect 21821 6267 21879 6273
rect 23109 6307 23167 6313
rect 23109 6273 23121 6307
rect 23155 6273 23167 6307
rect 23109 6267 23167 6273
rect 21836 6236 21864 6267
rect 22278 6236 22284 6248
rect 21836 6208 22284 6236
rect 22278 6196 22284 6208
rect 22336 6236 22342 6248
rect 23124 6236 23152 6267
rect 23382 6264 23388 6316
rect 23440 6304 23446 6316
rect 26206 6304 26234 6412
rect 38654 6400 38660 6412
rect 38712 6400 38718 6452
rect 23440 6276 26234 6304
rect 23440 6264 23446 6276
rect 22336 6208 23152 6236
rect 22336 6196 22342 6208
rect 1104 6010 48852 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 48852 6010
rect 1104 5936 48852 5958
rect 3418 5856 3424 5908
rect 3476 5896 3482 5908
rect 3476 5868 6914 5896
rect 3476 5856 3482 5868
rect 6886 5828 6914 5868
rect 23474 5856 23480 5908
rect 23532 5896 23538 5908
rect 24673 5899 24731 5905
rect 24673 5896 24685 5899
rect 23532 5868 24685 5896
rect 23532 5856 23538 5868
rect 24673 5865 24685 5868
rect 24719 5896 24731 5899
rect 25041 5899 25099 5905
rect 25041 5896 25053 5899
rect 24719 5868 25053 5896
rect 24719 5865 24731 5868
rect 24673 5859 24731 5865
rect 25041 5865 25053 5868
rect 25087 5865 25099 5899
rect 25041 5859 25099 5865
rect 25406 5856 25412 5908
rect 25464 5896 25470 5908
rect 25501 5899 25559 5905
rect 25501 5896 25513 5899
rect 25464 5868 25513 5896
rect 25464 5856 25470 5868
rect 25501 5865 25513 5868
rect 25547 5865 25559 5899
rect 25501 5859 25559 5865
rect 26970 5828 26976 5840
rect 6886 5800 26976 5828
rect 26970 5788 26976 5800
rect 27028 5788 27034 5840
rect 25225 5763 25283 5769
rect 25225 5729 25237 5763
rect 25271 5760 25283 5763
rect 48133 5763 48191 5769
rect 48133 5760 48145 5763
rect 25271 5732 48145 5760
rect 25271 5729 25283 5732
rect 25225 5723 25283 5729
rect 48133 5729 48145 5732
rect 48179 5729 48191 5763
rect 48133 5723 48191 5729
rect 2130 5652 2136 5704
rect 2188 5692 2194 5704
rect 2317 5695 2375 5701
rect 2317 5692 2329 5695
rect 2188 5664 2329 5692
rect 2188 5652 2194 5664
rect 2317 5661 2329 5664
rect 2363 5661 2375 5695
rect 2317 5655 2375 5661
rect 2961 5695 3019 5701
rect 2961 5661 2973 5695
rect 3007 5692 3019 5695
rect 25317 5695 25375 5701
rect 3007 5664 22094 5692
rect 3007 5661 3019 5664
rect 2961 5655 3019 5661
rect 3050 5556 3056 5568
rect 3011 5528 3056 5556
rect 3050 5516 3056 5528
rect 3108 5516 3114 5568
rect 22066 5556 22094 5664
rect 25317 5661 25329 5695
rect 25363 5692 25375 5695
rect 25866 5692 25872 5704
rect 25363 5664 25872 5692
rect 25363 5661 25375 5664
rect 25317 5655 25375 5661
rect 25866 5652 25872 5664
rect 25924 5652 25930 5704
rect 47394 5692 47400 5704
rect 47355 5664 47400 5692
rect 47394 5652 47400 5664
rect 47452 5652 47458 5704
rect 25041 5627 25099 5633
rect 25041 5593 25053 5627
rect 25087 5624 25099 5627
rect 35342 5624 35348 5636
rect 25087 5596 35348 5624
rect 25087 5593 25099 5596
rect 25041 5587 25099 5593
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 47946 5624 47952 5636
rect 47907 5596 47952 5624
rect 47946 5584 47952 5596
rect 48004 5584 48010 5636
rect 26786 5556 26792 5568
rect 22066 5528 26792 5556
rect 26786 5516 26792 5528
rect 26844 5516 26850 5568
rect 1104 5466 48852 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 48852 5466
rect 1104 5392 48852 5414
rect 2317 5287 2375 5293
rect 2317 5253 2329 5287
rect 2363 5284 2375 5287
rect 3050 5284 3056 5296
rect 2363 5256 3056 5284
rect 2363 5253 2375 5256
rect 2317 5247 2375 5253
rect 3050 5244 3056 5256
rect 3108 5244 3114 5296
rect 2130 5216 2136 5228
rect 2091 5188 2136 5216
rect 2130 5176 2136 5188
rect 2188 5176 2194 5228
rect 46842 5216 46848 5228
rect 46755 5188 46848 5216
rect 46842 5176 46848 5188
rect 46900 5216 46906 5228
rect 47486 5216 47492 5228
rect 46900 5188 47492 5216
rect 46900 5176 46906 5188
rect 47486 5176 47492 5188
rect 47544 5176 47550 5228
rect 47578 5176 47584 5228
rect 47636 5216 47642 5228
rect 48222 5216 48228 5228
rect 47636 5188 48228 5216
rect 47636 5176 47642 5188
rect 48222 5176 48228 5188
rect 48280 5176 48286 5228
rect 2774 5148 2780 5160
rect 2735 5120 2780 5148
rect 2774 5108 2780 5120
rect 2832 5108 2838 5160
rect 36354 5108 36360 5160
rect 36412 5148 36418 5160
rect 47026 5148 47032 5160
rect 36412 5120 47032 5148
rect 36412 5108 36418 5120
rect 47026 5108 47032 5120
rect 47084 5108 47090 5160
rect 1394 4972 1400 5024
rect 1452 5012 1458 5024
rect 1673 5015 1731 5021
rect 1673 5012 1685 5015
rect 1452 4984 1685 5012
rect 1452 4972 1458 4984
rect 1673 4981 1685 4984
rect 1719 4981 1731 5015
rect 46934 5012 46940 5024
rect 46895 4984 46940 5012
rect 1673 4975 1731 4981
rect 46934 4972 46940 4984
rect 46992 4972 46998 5024
rect 47670 5012 47676 5024
rect 47631 4984 47676 5012
rect 47670 4972 47676 4984
rect 47728 4972 47734 5024
rect 1104 4922 48852 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 48852 4922
rect 1104 4848 48852 4870
rect 35434 4768 35440 4820
rect 35492 4808 35498 4820
rect 45554 4808 45560 4820
rect 35492 4780 45560 4808
rect 35492 4768 35498 4780
rect 45554 4768 45560 4780
rect 45612 4768 45618 4820
rect 47394 4740 47400 4752
rect 46308 4712 47400 4740
rect 1394 4672 1400 4684
rect 1355 4644 1400 4672
rect 1394 4632 1400 4644
rect 1452 4632 1458 4684
rect 1581 4675 1639 4681
rect 1581 4641 1593 4675
rect 1627 4672 1639 4675
rect 3881 4675 3939 4681
rect 3881 4672 3893 4675
rect 1627 4644 3893 4672
rect 1627 4641 1639 4644
rect 1581 4635 1639 4641
rect 3881 4641 3893 4644
rect 3927 4641 3939 4675
rect 3881 4635 3939 4641
rect 21910 4632 21916 4684
rect 21968 4672 21974 4684
rect 22005 4675 22063 4681
rect 22005 4672 22017 4675
rect 21968 4644 22017 4672
rect 21968 4632 21974 4644
rect 22005 4641 22017 4644
rect 22051 4641 22063 4675
rect 22005 4635 22063 4641
rect 34790 4632 34796 4684
rect 34848 4672 34854 4684
rect 37366 4672 37372 4684
rect 34848 4644 37372 4672
rect 34848 4632 34854 4644
rect 37366 4632 37372 4644
rect 37424 4632 37430 4684
rect 41877 4675 41935 4681
rect 41877 4641 41889 4675
rect 41923 4672 41935 4675
rect 43070 4672 43076 4684
rect 41923 4644 43076 4672
rect 41923 4641 41935 4644
rect 41877 4635 41935 4641
rect 43070 4632 43076 4644
rect 43128 4632 43134 4684
rect 43254 4672 43260 4684
rect 43215 4644 43260 4672
rect 43254 4632 43260 4644
rect 43312 4632 43318 4684
rect 46308 4681 46336 4712
rect 47394 4700 47400 4712
rect 47452 4700 47458 4752
rect 46293 4675 46351 4681
rect 46293 4641 46305 4675
rect 46339 4641 46351 4675
rect 46293 4635 46351 4641
rect 46477 4675 46535 4681
rect 46477 4641 46489 4675
rect 46523 4672 46535 4675
rect 47670 4672 47676 4684
rect 46523 4644 47676 4672
rect 46523 4641 46535 4644
rect 46477 4635 46535 4641
rect 47670 4632 47676 4644
rect 47728 4632 47734 4684
rect 48130 4672 48136 4684
rect 48091 4644 48136 4672
rect 48130 4632 48136 4644
rect 48188 4632 48194 4684
rect 3234 4604 3240 4616
rect 3195 4576 3240 4604
rect 3234 4564 3240 4576
rect 3292 4564 3298 4616
rect 3786 4604 3792 4616
rect 3747 4576 3792 4604
rect 3786 4564 3792 4576
rect 3844 4564 3850 4616
rect 6270 4604 6276 4616
rect 6231 4576 6276 4604
rect 6270 4564 6276 4576
rect 6328 4564 6334 4616
rect 6917 4607 6975 4613
rect 6917 4573 6929 4607
rect 6963 4604 6975 4607
rect 7190 4604 7196 4616
rect 6963 4576 7196 4604
rect 6963 4573 6975 4576
rect 6917 4567 6975 4573
rect 7190 4564 7196 4576
rect 7248 4564 7254 4616
rect 8018 4604 8024 4616
rect 7979 4576 8024 4604
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 30466 4604 30472 4616
rect 30427 4576 30472 4604
rect 30466 4564 30472 4576
rect 30524 4564 30530 4616
rect 30834 4564 30840 4616
rect 30892 4604 30898 4616
rect 31113 4607 31171 4613
rect 31113 4604 31125 4607
rect 30892 4576 31125 4604
rect 30892 4564 30898 4576
rect 31113 4573 31125 4576
rect 31159 4573 31171 4607
rect 31113 4567 31171 4573
rect 44726 4564 44732 4616
rect 44784 4604 44790 4616
rect 45189 4607 45247 4613
rect 45189 4604 45201 4607
rect 44784 4576 45201 4604
rect 44784 4564 44790 4576
rect 45189 4573 45201 4576
rect 45235 4573 45247 4607
rect 45830 4604 45836 4616
rect 45791 4576 45836 4604
rect 45189 4567 45247 4573
rect 45830 4564 45836 4576
rect 45888 4564 45894 4616
rect 22186 4536 22192 4548
rect 22147 4508 22192 4536
rect 22186 4496 22192 4508
rect 22244 4496 22250 4548
rect 23845 4539 23903 4545
rect 23845 4505 23857 4539
rect 23891 4536 23903 4539
rect 34514 4536 34520 4548
rect 23891 4508 34520 4536
rect 23891 4505 23903 4508
rect 23845 4499 23903 4505
rect 34514 4496 34520 4508
rect 34572 4496 34578 4548
rect 42058 4536 42064 4548
rect 42019 4508 42064 4536
rect 42058 4496 42064 4508
rect 42116 4496 42122 4548
rect 8110 4468 8116 4480
rect 8071 4440 8116 4468
rect 8110 4428 8116 4440
rect 8168 4428 8174 4480
rect 1104 4378 48852 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 48852 4378
rect 1104 4304 48852 4326
rect 22186 4224 22192 4276
rect 22244 4264 22250 4276
rect 22649 4267 22707 4273
rect 22649 4264 22661 4267
rect 22244 4236 22661 4264
rect 22244 4224 22250 4236
rect 22649 4233 22661 4236
rect 22695 4233 22707 4267
rect 22649 4227 22707 4233
rect 42058 4224 42064 4276
rect 42116 4264 42122 4276
rect 42521 4267 42579 4273
rect 42521 4264 42533 4267
rect 42116 4236 42533 4264
rect 42116 4224 42122 4236
rect 42521 4233 42533 4236
rect 42567 4233 42579 4267
rect 42521 4227 42579 4233
rect 3418 4156 3424 4208
rect 3476 4196 3482 4208
rect 8110 4196 8116 4208
rect 3476 4168 6914 4196
rect 8071 4168 8116 4196
rect 3476 4156 3482 4168
rect 1946 4088 1952 4140
rect 2004 4128 2010 4140
rect 2041 4131 2099 4137
rect 2041 4128 2053 4131
rect 2004 4100 2053 4128
rect 2004 4088 2010 4100
rect 2041 4097 2053 4100
rect 2087 4097 2099 4131
rect 2682 4128 2688 4140
rect 2643 4100 2688 4128
rect 2041 4091 2099 4097
rect 2682 4088 2688 4100
rect 2740 4088 2746 4140
rect 6362 4128 6368 4140
rect 6323 4100 6368 4128
rect 6362 4088 6368 4100
rect 6420 4088 6426 4140
rect 2130 4020 2136 4072
rect 2188 4060 2194 4072
rect 6178 4060 6184 4072
rect 2188 4032 6184 4060
rect 2188 4020 2194 4032
rect 6178 4020 6184 4032
rect 6236 4020 6242 4072
rect 6886 4060 6914 4168
rect 8110 4156 8116 4168
rect 8168 4156 8174 4208
rect 10226 4156 10232 4208
rect 10284 4196 10290 4208
rect 17954 4196 17960 4208
rect 10284 4168 17960 4196
rect 10284 4156 10290 4168
rect 17954 4156 17960 4168
rect 18012 4156 18018 4208
rect 20548 4168 26234 4196
rect 7006 4088 7012 4140
rect 7064 4128 7070 4140
rect 7926 4128 7932 4140
rect 7064 4100 7109 4128
rect 7887 4100 7932 4128
rect 7064 4088 7070 4100
rect 7926 4088 7932 4100
rect 7984 4088 7990 4140
rect 11609 4131 11667 4137
rect 11609 4128 11621 4131
rect 9324 4100 11621 4128
rect 8389 4063 8447 4069
rect 8389 4060 8401 4063
rect 6886 4032 8401 4060
rect 8389 4029 8401 4032
rect 8435 4029 8447 4063
rect 8389 4023 8447 4029
rect 2498 3952 2504 4004
rect 2556 3992 2562 4004
rect 9324 3992 9352 4100
rect 11609 4097 11621 4100
rect 11655 4097 11667 4131
rect 12526 4128 12532 4140
rect 12487 4100 12532 4128
rect 11609 4091 11667 4097
rect 12526 4088 12532 4100
rect 12584 4088 12590 4140
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 20548 4128 20576 4168
rect 14976 4100 20576 4128
rect 14976 4088 14982 4100
rect 22554 4088 22560 4140
rect 22612 4128 22618 4140
rect 26206 4128 26234 4168
rect 29454 4156 29460 4208
rect 29512 4196 29518 4208
rect 29512 4168 30788 4196
rect 29512 4156 29518 4168
rect 30190 4128 30196 4140
rect 22612 4100 22657 4128
rect 26206 4100 30196 4128
rect 22612 4088 22618 4100
rect 30190 4088 30196 4100
rect 30248 4088 30254 4140
rect 30760 4137 30788 4168
rect 36280 4168 36492 4196
rect 30745 4131 30803 4137
rect 30745 4097 30757 4131
rect 30791 4128 30803 4131
rect 31294 4128 31300 4140
rect 30791 4100 31300 4128
rect 30791 4097 30803 4100
rect 30745 4091 30803 4097
rect 31294 4088 31300 4100
rect 31352 4088 31358 4140
rect 31389 4131 31447 4137
rect 31389 4097 31401 4131
rect 31435 4097 31447 4131
rect 36280 4128 36308 4168
rect 31389 4091 31447 4097
rect 35866 4100 36308 4128
rect 36357 4131 36415 4137
rect 10686 4060 10692 4072
rect 2556 3964 9352 3992
rect 9416 4032 10692 4060
rect 2556 3952 2562 3964
rect 1578 3924 1584 3936
rect 1539 3896 1584 3924
rect 1578 3884 1584 3896
rect 1636 3884 1642 3936
rect 1670 3884 1676 3936
rect 1728 3924 1734 3936
rect 2133 3927 2191 3933
rect 2133 3924 2145 3927
rect 1728 3896 2145 3924
rect 1728 3884 1734 3896
rect 2133 3893 2145 3896
rect 2179 3893 2191 3927
rect 2133 3887 2191 3893
rect 2777 3927 2835 3933
rect 2777 3893 2789 3927
rect 2823 3924 2835 3927
rect 2866 3924 2872 3936
rect 2823 3896 2872 3924
rect 2823 3893 2835 3896
rect 2777 3887 2835 3893
rect 2866 3884 2872 3896
rect 2924 3884 2930 3936
rect 3510 3884 3516 3936
rect 3568 3924 3574 3936
rect 3789 3927 3847 3933
rect 3789 3924 3801 3927
rect 3568 3896 3801 3924
rect 3568 3884 3574 3896
rect 3789 3893 3801 3896
rect 3835 3893 3847 3927
rect 3789 3887 3847 3893
rect 5166 3884 5172 3936
rect 5224 3924 5230 3936
rect 5445 3927 5503 3933
rect 5445 3924 5457 3927
rect 5224 3896 5457 3924
rect 5224 3884 5230 3896
rect 5445 3893 5457 3896
rect 5491 3893 5503 3927
rect 5445 3887 5503 3893
rect 5534 3884 5540 3936
rect 5592 3924 5598 3936
rect 6457 3927 6515 3933
rect 6457 3924 6469 3927
rect 5592 3896 6469 3924
rect 5592 3884 5598 3896
rect 6457 3893 6469 3896
rect 6503 3893 6515 3927
rect 7098 3924 7104 3936
rect 7059 3896 7104 3924
rect 6457 3887 6515 3893
rect 7098 3884 7104 3896
rect 7156 3884 7162 3936
rect 7926 3884 7932 3936
rect 7984 3924 7990 3936
rect 9416 3924 9444 4032
rect 10686 4020 10692 4032
rect 10744 4060 10750 4072
rect 12434 4060 12440 4072
rect 10744 4032 12440 4060
rect 10744 4020 10750 4032
rect 12434 4020 12440 4032
rect 12492 4020 12498 4072
rect 13170 4060 13176 4072
rect 13131 4032 13176 4060
rect 13170 4020 13176 4032
rect 13228 4020 13234 4072
rect 13357 4063 13415 4069
rect 13357 4029 13369 4063
rect 13403 4029 13415 4063
rect 13357 4023 13415 4029
rect 10318 3952 10324 4004
rect 10376 3992 10382 4004
rect 12342 3992 12348 4004
rect 10376 3964 12348 3992
rect 10376 3952 10382 3964
rect 12342 3952 12348 3964
rect 12400 3952 12406 4004
rect 12621 3995 12679 4001
rect 12621 3961 12633 3995
rect 12667 3992 12679 3995
rect 13372 3992 13400 4023
rect 13538 4020 13544 4072
rect 13596 4060 13602 4072
rect 13633 4063 13691 4069
rect 13633 4060 13645 4063
rect 13596 4032 13645 4060
rect 13596 4020 13602 4032
rect 13633 4029 13645 4032
rect 13679 4029 13691 4063
rect 13633 4023 13691 4029
rect 17218 4020 17224 4072
rect 17276 4060 17282 4072
rect 22462 4060 22468 4072
rect 17276 4032 22468 4060
rect 17276 4020 17282 4032
rect 22462 4020 22468 4032
rect 22520 4020 22526 4072
rect 26418 4060 26424 4072
rect 22572 4032 26424 4060
rect 22572 3992 22600 4032
rect 26418 4020 26424 4032
rect 26476 4020 26482 4072
rect 28350 4020 28356 4072
rect 28408 4060 28414 4072
rect 31404 4060 31432 4091
rect 28408 4032 31432 4060
rect 28408 4020 28414 4032
rect 12667 3964 13400 3992
rect 15948 3964 22600 3992
rect 12667 3961 12679 3964
rect 12621 3955 12679 3961
rect 7984 3896 9444 3924
rect 11701 3927 11759 3933
rect 7984 3884 7990 3896
rect 11701 3893 11713 3927
rect 11747 3924 11759 3927
rect 11882 3924 11888 3936
rect 11747 3896 11888 3924
rect 11747 3893 11759 3896
rect 11701 3887 11759 3893
rect 11882 3884 11888 3896
rect 11940 3884 11946 3936
rect 12526 3884 12532 3936
rect 12584 3924 12590 3936
rect 15948 3924 15976 3964
rect 24394 3952 24400 4004
rect 24452 3992 24458 4004
rect 35866 3992 35894 4100
rect 36357 4097 36369 4131
rect 36403 4097 36415 4131
rect 36464 4128 36492 4168
rect 43364 4168 43576 4196
rect 37826 4128 37832 4140
rect 36464 4100 37832 4128
rect 36357 4091 36415 4097
rect 36372 4060 36400 4091
rect 37826 4088 37832 4100
rect 37884 4088 37890 4140
rect 40957 4131 41015 4137
rect 40957 4097 40969 4131
rect 41003 4128 41015 4131
rect 42334 4128 42340 4140
rect 41003 4100 42340 4128
rect 41003 4097 41015 4100
rect 40957 4091 41015 4097
rect 42334 4088 42340 4100
rect 42392 4088 42398 4140
rect 42426 4088 42432 4140
rect 42484 4128 42490 4140
rect 42484 4100 42529 4128
rect 42484 4088 42490 4100
rect 43364 4060 43392 4168
rect 43441 4131 43499 4137
rect 43441 4097 43453 4131
rect 43487 4097 43499 4131
rect 43548 4128 43576 4168
rect 46750 4156 46756 4208
rect 46808 4196 46814 4208
rect 47949 4199 48007 4205
rect 47949 4196 47961 4199
rect 46808 4168 47961 4196
rect 46808 4156 46814 4168
rect 47949 4165 47961 4168
rect 47995 4165 48007 4199
rect 47949 4159 48007 4165
rect 43990 4128 43996 4140
rect 43548 4100 43996 4128
rect 43441 4091 43499 4097
rect 36372 4032 43392 4060
rect 24452 3964 35894 3992
rect 24452 3952 24458 3964
rect 12584 3896 15976 3924
rect 12584 3884 12590 3896
rect 17310 3884 17316 3936
rect 17368 3924 17374 3936
rect 17589 3927 17647 3933
rect 17589 3924 17601 3927
rect 17368 3896 17601 3924
rect 17368 3884 17374 3896
rect 17589 3893 17601 3896
rect 17635 3893 17647 3927
rect 20990 3924 20996 3936
rect 20951 3896 20996 3924
rect 17589 3887 17647 3893
rect 20990 3884 20996 3896
rect 21048 3884 21054 3936
rect 23382 3884 23388 3936
rect 23440 3924 23446 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23440 3896 23673 3924
rect 23440 3884 23446 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 25682 3884 25688 3936
rect 25740 3924 25746 3936
rect 25961 3927 26019 3933
rect 25961 3924 25973 3927
rect 25740 3896 25973 3924
rect 25740 3884 25746 3896
rect 25961 3893 25973 3896
rect 26007 3893 26019 3927
rect 25961 3887 26019 3893
rect 29730 3884 29736 3936
rect 29788 3924 29794 3936
rect 30009 3927 30067 3933
rect 30009 3924 30021 3927
rect 29788 3896 30021 3924
rect 29788 3884 29794 3896
rect 30009 3893 30021 3896
rect 30055 3893 30067 3927
rect 30009 3887 30067 3893
rect 30837 3927 30895 3933
rect 30837 3893 30849 3927
rect 30883 3924 30895 3927
rect 31018 3924 31024 3936
rect 30883 3896 31024 3924
rect 30883 3893 30895 3896
rect 30837 3887 30895 3893
rect 31018 3884 31024 3896
rect 31076 3884 31082 3936
rect 31478 3924 31484 3936
rect 31439 3896 31484 3924
rect 31478 3884 31484 3896
rect 31536 3884 31542 3936
rect 32122 3884 32128 3936
rect 32180 3924 32186 3936
rect 32401 3927 32459 3933
rect 32401 3924 32413 3927
rect 32180 3896 32413 3924
rect 32180 3884 32186 3896
rect 32401 3893 32413 3896
rect 32447 3893 32459 3927
rect 32401 3887 32459 3893
rect 36262 3884 36268 3936
rect 36320 3924 36326 3936
rect 36449 3927 36507 3933
rect 36449 3924 36461 3927
rect 36320 3896 36461 3924
rect 36320 3884 36326 3896
rect 36449 3893 36461 3896
rect 36495 3893 36507 3927
rect 36449 3887 36507 3893
rect 37921 3927 37979 3933
rect 37921 3893 37933 3927
rect 37967 3924 37979 3927
rect 38746 3924 38752 3936
rect 37967 3896 38752 3924
rect 37967 3893 37979 3896
rect 37921 3887 37979 3893
rect 38746 3884 38752 3896
rect 38804 3884 38810 3936
rect 40770 3884 40776 3936
rect 40828 3924 40834 3936
rect 41049 3927 41107 3933
rect 41049 3924 41061 3927
rect 40828 3896 41061 3924
rect 40828 3884 40834 3896
rect 41049 3893 41061 3896
rect 41095 3893 41107 3927
rect 41049 3887 41107 3893
rect 41785 3927 41843 3933
rect 41785 3893 41797 3927
rect 41831 3924 41843 3927
rect 42426 3924 42432 3936
rect 41831 3896 42432 3924
rect 41831 3893 41843 3896
rect 41785 3887 41843 3893
rect 42426 3884 42432 3896
rect 42484 3884 42490 3936
rect 43456 3924 43484 4091
rect 43990 4088 43996 4100
rect 44048 4088 44054 4140
rect 45462 4088 45468 4140
rect 45520 4128 45526 4140
rect 46385 4131 46443 4137
rect 46385 4128 46397 4131
rect 45520 4100 46397 4128
rect 45520 4088 45526 4100
rect 46385 4097 46397 4100
rect 46431 4097 46443 4131
rect 46385 4091 46443 4097
rect 43806 4020 43812 4072
rect 43864 4060 43870 4072
rect 44085 4063 44143 4069
rect 44085 4060 44097 4063
rect 43864 4032 44097 4060
rect 43864 4020 43870 4032
rect 44085 4029 44097 4032
rect 44131 4029 44143 4063
rect 44085 4023 44143 4029
rect 44269 4063 44327 4069
rect 44269 4029 44281 4063
rect 44315 4029 44327 4063
rect 44269 4023 44327 4029
rect 43533 3995 43591 4001
rect 43533 3961 43545 3995
rect 43579 3992 43591 3995
rect 44284 3992 44312 4023
rect 44450 4020 44456 4072
rect 44508 4060 44514 4072
rect 44545 4063 44603 4069
rect 44545 4060 44557 4063
rect 44508 4032 44557 4060
rect 44508 4020 44514 4032
rect 44545 4029 44557 4032
rect 44591 4029 44603 4063
rect 44545 4023 44603 4029
rect 43579 3964 44312 3992
rect 43579 3961 43591 3964
rect 43533 3955 43591 3961
rect 44818 3952 44824 4004
rect 44876 3992 44882 4004
rect 46842 3992 46848 4004
rect 44876 3964 46848 3992
rect 44876 3952 44882 3964
rect 46842 3952 46848 3964
rect 46900 3952 46906 4004
rect 45738 3924 45744 3936
rect 43456 3896 45744 3924
rect 45738 3884 45744 3896
rect 45796 3884 45802 3936
rect 46198 3884 46204 3936
rect 46256 3924 46262 3936
rect 46477 3927 46535 3933
rect 46477 3924 46489 3927
rect 46256 3896 46489 3924
rect 46256 3884 46262 3896
rect 46477 3893 46489 3896
rect 46523 3893 46535 3927
rect 48038 3924 48044 3936
rect 47999 3896 48044 3924
rect 46477 3887 46535 3893
rect 48038 3884 48044 3896
rect 48096 3884 48102 3936
rect 1104 3834 48852 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 48852 3834
rect 1104 3760 48852 3782
rect 2958 3680 2964 3732
rect 3016 3720 3022 3732
rect 12434 3720 12440 3732
rect 3016 3692 12440 3720
rect 3016 3680 3022 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 17218 3720 17224 3732
rect 12544 3692 17224 3720
rect 7926 3652 7932 3664
rect 4356 3624 7932 3652
rect 1581 3587 1639 3593
rect 1581 3553 1593 3587
rect 1627 3584 1639 3587
rect 1670 3584 1676 3596
rect 1627 3556 1676 3584
rect 1627 3553 1639 3556
rect 1581 3547 1639 3553
rect 1670 3544 1676 3556
rect 1728 3544 1734 3596
rect 1854 3584 1860 3596
rect 1815 3556 1860 3584
rect 1854 3544 1860 3556
rect 1912 3544 1918 3596
rect 1397 3519 1455 3525
rect 1397 3485 1409 3519
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 1412 3448 1440 3479
rect 3878 3476 3884 3528
rect 3936 3516 3942 3528
rect 4356 3525 4384 3624
rect 7926 3612 7932 3624
rect 7984 3612 7990 3664
rect 8018 3612 8024 3664
rect 8076 3652 8082 3664
rect 12544 3652 12572 3692
rect 17218 3680 17224 3692
rect 17276 3680 17282 3732
rect 17586 3680 17592 3732
rect 17644 3720 17650 3732
rect 19426 3720 19432 3732
rect 17644 3692 19432 3720
rect 17644 3680 17650 3692
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 22646 3720 22652 3732
rect 22607 3692 22652 3720
rect 22646 3680 22652 3692
rect 22704 3680 22710 3732
rect 23290 3680 23296 3732
rect 23348 3720 23354 3732
rect 33778 3720 33784 3732
rect 23348 3692 33784 3720
rect 23348 3680 23354 3692
rect 33778 3680 33784 3692
rect 33836 3680 33842 3732
rect 43070 3720 43076 3732
rect 43031 3692 43076 3720
rect 43070 3680 43076 3692
rect 43128 3680 43134 3732
rect 43806 3720 43812 3732
rect 43767 3692 43812 3720
rect 43806 3680 43812 3692
rect 43864 3680 43870 3732
rect 43990 3680 43996 3732
rect 44048 3720 44054 3732
rect 47578 3720 47584 3732
rect 44048 3692 47584 3720
rect 44048 3680 44054 3692
rect 47578 3680 47584 3692
rect 47636 3680 47642 3732
rect 30006 3652 30012 3664
rect 8076 3624 12572 3652
rect 12728 3624 18460 3652
rect 8076 3612 8082 3624
rect 5166 3584 5172 3596
rect 5127 3556 5172 3584
rect 5166 3544 5172 3556
rect 5224 3544 5230 3596
rect 5353 3587 5411 3593
rect 5353 3553 5365 3587
rect 5399 3584 5411 3587
rect 5534 3584 5540 3596
rect 5399 3556 5540 3584
rect 5399 3553 5411 3556
rect 5353 3547 5411 3553
rect 5534 3544 5540 3556
rect 5592 3544 5598 3596
rect 6549 3587 6607 3593
rect 6549 3553 6561 3587
rect 6595 3553 6607 3587
rect 6549 3547 6607 3553
rect 4341 3519 4399 3525
rect 3936 3488 4108 3516
rect 3936 3476 3942 3488
rect 3970 3448 3976 3460
rect 1412 3420 3976 3448
rect 3970 3408 3976 3420
rect 4028 3408 4034 3460
rect 4080 3448 4108 3488
rect 4341 3485 4353 3519
rect 4387 3485 4399 3519
rect 4341 3479 4399 3485
rect 4080 3420 4568 3448
rect 3694 3340 3700 3392
rect 3752 3380 3758 3392
rect 4433 3383 4491 3389
rect 4433 3380 4445 3383
rect 3752 3352 4445 3380
rect 3752 3340 3758 3352
rect 4433 3349 4445 3352
rect 4479 3349 4491 3383
rect 4540 3380 4568 3420
rect 5166 3408 5172 3460
rect 5224 3448 5230 3460
rect 6564 3448 6592 3547
rect 7006 3544 7012 3596
rect 7064 3584 7070 3596
rect 12728 3584 12756 3624
rect 7064 3556 12756 3584
rect 7064 3544 7070 3556
rect 7484 3525 7512 3556
rect 12802 3544 12808 3596
rect 12860 3584 12866 3596
rect 18322 3584 18328 3596
rect 12860 3556 12905 3584
rect 13096 3556 18328 3584
rect 12860 3544 12866 3556
rect 7469 3519 7527 3525
rect 7469 3485 7481 3519
rect 7515 3485 7527 3519
rect 7469 3479 7527 3485
rect 9030 3476 9036 3528
rect 9088 3516 9094 3528
rect 10502 3516 10508 3528
rect 9088 3488 10508 3516
rect 9088 3476 9094 3488
rect 10502 3476 10508 3488
rect 10560 3476 10566 3528
rect 11698 3516 11704 3528
rect 11659 3488 11704 3516
rect 11698 3476 11704 3488
rect 11756 3476 11762 3528
rect 5224 3420 6592 3448
rect 5224 3408 5230 3420
rect 6914 3408 6920 3460
rect 6972 3448 6978 3460
rect 7561 3451 7619 3457
rect 7561 3448 7573 3451
rect 6972 3420 7573 3448
rect 6972 3408 6978 3420
rect 7561 3417 7573 3420
rect 7607 3417 7619 3451
rect 7561 3411 7619 3417
rect 11882 3408 11888 3460
rect 11940 3448 11946 3460
rect 11940 3420 11985 3448
rect 11940 3408 11946 3420
rect 12434 3408 12440 3460
rect 12492 3448 12498 3460
rect 13096 3448 13124 3556
rect 18322 3544 18328 3556
rect 18380 3544 18386 3596
rect 14461 3519 14519 3525
rect 14461 3485 14473 3519
rect 14507 3516 14519 3519
rect 14918 3516 14924 3528
rect 14507 3488 14924 3516
rect 14507 3485 14519 3488
rect 14461 3479 14519 3485
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 15102 3516 15108 3528
rect 15063 3488 15108 3516
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 17681 3519 17739 3525
rect 16960 3516 17080 3518
rect 17681 3516 17693 3519
rect 16500 3490 17693 3516
rect 16500 3488 16988 3490
rect 17052 3488 17693 3490
rect 12492 3420 13124 3448
rect 14553 3451 14611 3457
rect 12492 3408 12498 3420
rect 14553 3417 14565 3451
rect 14599 3448 14611 3451
rect 15289 3451 15347 3457
rect 15289 3448 15301 3451
rect 14599 3420 15301 3448
rect 14599 3417 14611 3420
rect 14553 3411 14611 3417
rect 15289 3417 15301 3420
rect 15335 3417 15347 3451
rect 16500 3448 16528 3488
rect 17681 3485 17693 3488
rect 17727 3485 17739 3519
rect 17681 3479 17739 3485
rect 15289 3411 15347 3417
rect 15396 3420 16528 3448
rect 16945 3451 17003 3457
rect 11514 3380 11520 3392
rect 4540 3352 11520 3380
rect 4433 3343 4491 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 11606 3340 11612 3392
rect 11664 3380 11670 3392
rect 15396 3380 15424 3420
rect 16945 3417 16957 3451
rect 16991 3417 17003 3451
rect 16945 3411 17003 3417
rect 11664 3352 15424 3380
rect 11664 3340 11670 3352
rect 15470 3340 15476 3392
rect 15528 3380 15534 3392
rect 16960 3380 16988 3411
rect 15528 3352 16988 3380
rect 15528 3340 15534 3352
rect 17494 3340 17500 3392
rect 17552 3380 17558 3392
rect 17773 3383 17831 3389
rect 17773 3380 17785 3383
rect 17552 3352 17785 3380
rect 17552 3340 17558 3352
rect 17773 3349 17785 3352
rect 17819 3349 17831 3383
rect 18432 3380 18460 3624
rect 19628 3624 30012 3652
rect 19628 3525 19656 3624
rect 30006 3612 30012 3624
rect 30064 3612 30070 3664
rect 30190 3612 30196 3664
rect 30248 3652 30254 3664
rect 32398 3652 32404 3664
rect 30248 3624 32404 3652
rect 30248 3612 30254 3624
rect 32398 3612 32404 3624
rect 32456 3612 32462 3664
rect 35802 3612 35808 3664
rect 35860 3652 35866 3664
rect 45462 3652 45468 3664
rect 35860 3624 45468 3652
rect 35860 3612 35866 3624
rect 45462 3612 45468 3624
rect 45520 3612 45526 3664
rect 20622 3544 20628 3596
rect 20680 3584 20686 3596
rect 20717 3587 20775 3593
rect 20717 3584 20729 3587
rect 20680 3556 20729 3584
rect 20680 3544 20686 3556
rect 20717 3553 20729 3556
rect 20763 3553 20775 3587
rect 20717 3547 20775 3553
rect 22462 3544 22468 3596
rect 22520 3584 22526 3596
rect 25498 3584 25504 3596
rect 22520 3556 25504 3584
rect 22520 3544 22526 3556
rect 25498 3544 25504 3556
rect 25556 3544 25562 3596
rect 25682 3584 25688 3596
rect 25643 3556 25688 3584
rect 25682 3544 25688 3556
rect 25740 3544 25746 3596
rect 26418 3584 26424 3596
rect 26379 3556 26424 3584
rect 26418 3544 26424 3556
rect 26476 3544 26482 3596
rect 30834 3584 30840 3596
rect 29564 3556 30512 3584
rect 30795 3556 30840 3584
rect 29564 3528 29592 3556
rect 19613 3519 19671 3525
rect 19613 3485 19625 3519
rect 19659 3485 19671 3519
rect 20254 3516 20260 3528
rect 20215 3488 20260 3516
rect 19613 3479 19671 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 22833 3519 22891 3525
rect 22833 3485 22845 3519
rect 22879 3516 22891 3519
rect 23198 3516 23204 3528
rect 22879 3488 23204 3516
rect 22879 3485 22891 3488
rect 22833 3479 22891 3485
rect 23198 3476 23204 3488
rect 23256 3476 23262 3528
rect 23290 3476 23296 3528
rect 23348 3516 23354 3528
rect 29546 3516 29552 3528
rect 23348 3488 23393 3516
rect 29507 3488 29552 3516
rect 23348 3476 23354 3488
rect 29546 3476 29552 3488
rect 29604 3476 29610 3528
rect 30190 3516 30196 3528
rect 30151 3488 30196 3516
rect 30190 3476 30196 3488
rect 30248 3476 30254 3528
rect 19705 3451 19763 3457
rect 19705 3417 19717 3451
rect 19751 3448 19763 3451
rect 20441 3451 20499 3457
rect 20441 3448 20453 3451
rect 19751 3420 20453 3448
rect 19751 3417 19763 3420
rect 19705 3411 19763 3417
rect 20441 3417 20453 3420
rect 20487 3417 20499 3451
rect 25869 3451 25927 3457
rect 20441 3411 20499 3417
rect 22066 3420 23704 3448
rect 22066 3380 22094 3420
rect 18432 3352 22094 3380
rect 23385 3383 23443 3389
rect 17773 3343 17831 3349
rect 23385 3349 23397 3383
rect 23431 3380 23443 3383
rect 23566 3380 23572 3392
rect 23431 3352 23572 3380
rect 23431 3349 23443 3352
rect 23385 3343 23443 3349
rect 23566 3340 23572 3352
rect 23624 3340 23630 3392
rect 23676 3380 23704 3420
rect 25869 3417 25881 3451
rect 25915 3448 25927 3451
rect 26142 3448 26148 3460
rect 25915 3420 26148 3448
rect 25915 3417 25927 3420
rect 25869 3411 25927 3417
rect 26142 3408 26148 3420
rect 26200 3408 26206 3460
rect 30484 3448 30512 3556
rect 30834 3544 30840 3556
rect 30892 3544 30898 3596
rect 31018 3584 31024 3596
rect 30979 3556 31024 3584
rect 31018 3544 31024 3556
rect 31076 3544 31082 3596
rect 31570 3584 31576 3596
rect 31531 3556 31576 3584
rect 31570 3544 31576 3556
rect 31628 3544 31634 3596
rect 36262 3584 36268 3596
rect 36223 3556 36268 3584
rect 36262 3544 36268 3556
rect 36320 3544 36326 3596
rect 36722 3584 36728 3596
rect 36683 3556 36728 3584
rect 36722 3544 36728 3556
rect 36780 3544 36786 3596
rect 40770 3584 40776 3596
rect 40731 3556 40776 3584
rect 40770 3544 40776 3556
rect 40828 3544 40834 3596
rect 41230 3584 41236 3596
rect 41191 3556 41236 3584
rect 41230 3544 41236 3556
rect 41288 3544 41294 3596
rect 44453 3587 44511 3593
rect 44453 3553 44465 3587
rect 44499 3584 44511 3587
rect 46017 3587 46075 3593
rect 46017 3584 46029 3587
rect 44499 3556 46029 3584
rect 44499 3553 44511 3556
rect 44453 3547 44511 3553
rect 46017 3553 46029 3556
rect 46063 3553 46075 3587
rect 46198 3584 46204 3596
rect 46159 3556 46204 3584
rect 46017 3547 46075 3553
rect 46198 3544 46204 3556
rect 46256 3544 46262 3596
rect 46382 3544 46388 3596
rect 46440 3584 46446 3596
rect 46477 3587 46535 3593
rect 46477 3584 46489 3587
rect 46440 3556 46489 3584
rect 46440 3544 46446 3556
rect 46477 3553 46489 3556
rect 46523 3553 46535 3587
rect 46477 3547 46535 3553
rect 36078 3516 36084 3528
rect 36039 3488 36084 3516
rect 36078 3476 36084 3488
rect 36136 3476 36142 3528
rect 38562 3476 38568 3528
rect 38620 3516 38626 3528
rect 38749 3519 38807 3525
rect 38749 3516 38761 3519
rect 38620 3488 38761 3516
rect 38620 3476 38626 3488
rect 38749 3485 38761 3488
rect 38795 3485 38807 3519
rect 38749 3479 38807 3485
rect 39945 3519 40003 3525
rect 39945 3485 39957 3519
rect 39991 3516 40003 3519
rect 40589 3519 40647 3525
rect 40589 3516 40601 3519
rect 39991 3488 40601 3516
rect 39991 3485 40003 3488
rect 39945 3479 40003 3485
rect 40589 3485 40601 3488
rect 40635 3485 40647 3519
rect 40589 3479 40647 3485
rect 45005 3519 45063 3525
rect 45005 3485 45017 3519
rect 45051 3485 45063 3519
rect 45005 3479 45063 3485
rect 33962 3448 33968 3460
rect 26896 3420 30420 3448
rect 30484 3420 33968 3448
rect 26896 3380 26924 3420
rect 23676 3352 26924 3380
rect 29641 3383 29699 3389
rect 29641 3349 29653 3383
rect 29687 3380 29699 3383
rect 29914 3380 29920 3392
rect 29687 3352 29920 3380
rect 29687 3349 29699 3352
rect 29641 3343 29699 3349
rect 29914 3340 29920 3352
rect 29972 3340 29978 3392
rect 30282 3380 30288 3392
rect 30243 3352 30288 3380
rect 30282 3340 30288 3352
rect 30340 3340 30346 3392
rect 30392 3380 30420 3420
rect 33962 3408 33968 3420
rect 34020 3408 34026 3460
rect 44818 3448 44824 3460
rect 35866 3420 44824 3448
rect 35866 3380 35894 3420
rect 44818 3408 44824 3420
rect 44876 3408 44882 3460
rect 45020 3448 45048 3479
rect 47210 3448 47216 3460
rect 45020 3420 47216 3448
rect 47210 3408 47216 3420
rect 47268 3408 47274 3460
rect 30392 3352 35894 3380
rect 42518 3340 42524 3392
rect 42576 3380 42582 3392
rect 43254 3380 43260 3392
rect 42576 3352 43260 3380
rect 42576 3340 42582 3352
rect 43254 3340 43260 3352
rect 43312 3340 43318 3392
rect 44910 3340 44916 3392
rect 44968 3380 44974 3392
rect 45097 3383 45155 3389
rect 45097 3380 45109 3383
rect 44968 3352 45109 3380
rect 44968 3340 44974 3352
rect 45097 3349 45109 3352
rect 45143 3349 45155 3383
rect 45097 3343 45155 3349
rect 1104 3290 48852 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 48852 3290
rect 1104 3216 48852 3238
rect 1949 3179 2007 3185
rect 1949 3145 1961 3179
rect 1995 3176 2007 3179
rect 2130 3176 2136 3188
rect 1995 3148 2136 3176
rect 1995 3145 2007 3148
rect 1949 3139 2007 3145
rect 2130 3136 2136 3148
rect 2188 3136 2194 3188
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 4798 3176 4804 3188
rect 2648 3148 4804 3176
rect 2648 3136 2654 3148
rect 4798 3136 4804 3148
rect 4856 3136 4862 3188
rect 11606 3176 11612 3188
rect 4908 3148 11612 3176
rect 1857 3111 1915 3117
rect 1857 3077 1869 3111
rect 1903 3108 1915 3111
rect 2774 3108 2780 3120
rect 1903 3080 2780 3108
rect 1903 3077 1915 3080
rect 1857 3071 1915 3077
rect 2774 3068 2780 3080
rect 2832 3068 2838 3120
rect 3694 3108 3700 3120
rect 3655 3080 3700 3108
rect 3694 3068 3700 3080
rect 3752 3068 3758 3120
rect 1946 3000 1952 3052
rect 2004 3040 2010 3052
rect 2593 3043 2651 3049
rect 2593 3040 2605 3043
rect 2004 3012 2605 3040
rect 2004 3000 2010 3012
rect 2593 3009 2605 3012
rect 2639 3009 2651 3043
rect 3510 3040 3516 3052
rect 3471 3012 3516 3040
rect 2593 3003 2651 3009
rect 3510 3000 3516 3012
rect 3568 3000 3574 3052
rect 2777 2975 2835 2981
rect 2777 2941 2789 2975
rect 2823 2972 2835 2975
rect 2958 2972 2964 2984
rect 2823 2944 2964 2972
rect 2823 2941 2835 2944
rect 2777 2935 2835 2941
rect 2958 2932 2964 2944
rect 3016 2932 3022 2984
rect 3234 2932 3240 2984
rect 3292 2972 3298 2984
rect 3973 2975 4031 2981
rect 3973 2972 3985 2975
rect 3292 2944 3985 2972
rect 3292 2932 3298 2944
rect 3973 2941 3985 2944
rect 4019 2941 4031 2975
rect 3973 2935 4031 2941
rect 658 2864 664 2916
rect 716 2904 722 2916
rect 716 2876 2084 2904
rect 716 2864 722 2876
rect 2056 2836 2084 2876
rect 2682 2864 2688 2916
rect 2740 2904 2746 2916
rect 4908 2904 4936 3148
rect 11606 3136 11612 3148
rect 11664 3136 11670 3188
rect 26694 3176 26700 3188
rect 11716 3148 26700 3176
rect 11716 3108 11744 3148
rect 26694 3136 26700 3148
rect 26752 3136 26758 3188
rect 30006 3136 30012 3188
rect 30064 3176 30070 3188
rect 30064 3148 32444 3176
rect 30064 3136 30070 3148
rect 16482 3108 16488 3120
rect 2740 2876 4936 2904
rect 5000 3080 11744 3108
rect 12268 3080 16488 3108
rect 2740 2864 2746 2876
rect 5000 2836 5028 3080
rect 6270 3000 6276 3052
rect 6328 3040 6334 3052
rect 6365 3043 6423 3049
rect 6365 3040 6377 3043
rect 6328 3012 6377 3040
rect 6328 3000 6334 3012
rect 6365 3009 6377 3012
rect 6411 3009 6423 3043
rect 6365 3003 6423 3009
rect 9674 3000 9680 3052
rect 9732 3040 9738 3052
rect 10045 3043 10103 3049
rect 10045 3040 10057 3043
rect 9732 3012 10057 3040
rect 9732 3000 9738 3012
rect 10045 3009 10057 3012
rect 10091 3009 10103 3043
rect 10226 3040 10232 3052
rect 10187 3012 10232 3040
rect 10045 3003 10103 3009
rect 10226 3000 10232 3012
rect 10284 3000 10290 3052
rect 11698 3000 11704 3052
rect 11756 3040 11762 3052
rect 11977 3043 12035 3049
rect 11977 3040 11989 3043
rect 11756 3012 11989 3040
rect 11756 3000 11762 3012
rect 11977 3009 11989 3012
rect 12023 3009 12035 3043
rect 11977 3003 12035 3009
rect 6549 2975 6607 2981
rect 6549 2941 6561 2975
rect 6595 2941 6607 2975
rect 6549 2935 6607 2941
rect 6564 2904 6592 2935
rect 6638 2932 6644 2984
rect 6696 2972 6702 2984
rect 6825 2975 6883 2981
rect 6825 2972 6837 2975
rect 6696 2944 6837 2972
rect 6696 2932 6702 2944
rect 6825 2941 6837 2944
rect 6871 2941 6883 2975
rect 6825 2935 6883 2941
rect 7742 2932 7748 2984
rect 7800 2972 7806 2984
rect 8665 2975 8723 2981
rect 8665 2972 8677 2975
rect 7800 2944 8677 2972
rect 7800 2932 7806 2944
rect 8665 2941 8677 2944
rect 8711 2941 8723 2975
rect 8665 2935 8723 2941
rect 8941 2975 8999 2981
rect 8941 2941 8953 2975
rect 8987 2972 8999 2975
rect 12268 2972 12296 3080
rect 16482 3068 16488 3080
rect 16540 3068 16546 3120
rect 17494 3108 17500 3120
rect 17455 3080 17500 3108
rect 17494 3068 17500 3080
rect 17552 3068 17558 3120
rect 17678 3068 17684 3120
rect 17736 3108 17742 3120
rect 23290 3108 23296 3120
rect 17736 3080 23296 3108
rect 17736 3068 17742 3080
rect 23290 3068 23296 3080
rect 23348 3068 23354 3120
rect 23566 3108 23572 3120
rect 23527 3080 23572 3108
rect 23566 3068 23572 3080
rect 23624 3068 23630 3120
rect 25498 3068 25504 3120
rect 25556 3108 25562 3120
rect 29454 3108 29460 3120
rect 25556 3080 29460 3108
rect 25556 3068 25562 3080
rect 29454 3068 29460 3080
rect 29512 3068 29518 3120
rect 29914 3068 29920 3120
rect 29972 3108 29978 3120
rect 29972 3080 30014 3108
rect 29972 3068 29978 3080
rect 31478 3068 31484 3120
rect 31536 3108 31542 3120
rect 32309 3111 32367 3117
rect 32309 3108 32321 3111
rect 31536 3080 32321 3108
rect 31536 3068 31542 3080
rect 32309 3077 32321 3080
rect 32355 3077 32367 3111
rect 32416 3108 32444 3148
rect 34238 3136 34244 3188
rect 34296 3176 34302 3188
rect 48038 3176 48044 3188
rect 34296 3148 48044 3176
rect 34296 3136 34302 3148
rect 48038 3136 48044 3148
rect 48096 3136 48102 3188
rect 34330 3108 34336 3120
rect 32416 3080 34336 3108
rect 32309 3071 32367 3077
rect 34330 3068 34336 3080
rect 34388 3108 34394 3120
rect 44910 3108 44916 3120
rect 34388 3080 41414 3108
rect 44871 3080 44916 3108
rect 34388 3068 34394 3080
rect 15102 3000 15108 3052
rect 15160 3040 15166 3052
rect 15289 3043 15347 3049
rect 15289 3040 15301 3043
rect 15160 3012 15301 3040
rect 15160 3000 15166 3012
rect 15289 3009 15301 3012
rect 15335 3009 15347 3043
rect 17310 3040 17316 3052
rect 17271 3012 17316 3040
rect 15289 3003 15347 3009
rect 17310 3000 17316 3012
rect 17368 3000 17374 3052
rect 20254 3000 20260 3052
rect 20312 3040 20318 3052
rect 20441 3043 20499 3049
rect 20441 3040 20453 3043
rect 20312 3012 20453 3040
rect 20312 3000 20318 3012
rect 20441 3009 20453 3012
rect 20487 3009 20499 3043
rect 20441 3003 20499 3009
rect 22554 3000 22560 3052
rect 22612 3040 22618 3052
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22612 3012 22753 3040
rect 22612 3000 22618 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 23382 3040 23388 3052
rect 23343 3012 23388 3040
rect 22741 3003 22799 3009
rect 23382 3000 23388 3012
rect 23440 3000 23446 3052
rect 26053 3043 26111 3049
rect 26053 3009 26065 3043
rect 26099 3040 26111 3043
rect 29546 3040 29552 3052
rect 26099 3012 29552 3040
rect 26099 3009 26111 3012
rect 26053 3003 26111 3009
rect 29546 3000 29552 3012
rect 29604 3000 29610 3052
rect 29730 3040 29736 3052
rect 29691 3012 29736 3040
rect 29730 3000 29736 3012
rect 29788 3000 29794 3052
rect 32122 3040 32128 3052
rect 32083 3012 32128 3040
rect 32122 3000 32128 3012
rect 32180 3000 32186 3052
rect 36078 3000 36084 3052
rect 36136 3040 36142 3052
rect 36265 3043 36323 3049
rect 36265 3040 36277 3043
rect 36136 3012 36277 3040
rect 36136 3000 36142 3012
rect 36265 3009 36277 3012
rect 36311 3009 36323 3043
rect 38562 3040 38568 3052
rect 38523 3012 38568 3040
rect 36265 3003 36323 3009
rect 38562 3000 38568 3012
rect 38620 3000 38626 3052
rect 41386 3040 41414 3080
rect 44910 3068 44916 3080
rect 44968 3068 44974 3120
rect 41509 3043 41567 3049
rect 41509 3040 41521 3043
rect 41386 3012 41521 3040
rect 41509 3009 41521 3012
rect 41555 3009 41567 3043
rect 42426 3040 42432 3052
rect 42387 3012 42432 3040
rect 41509 3003 41567 3009
rect 42426 3000 42432 3012
rect 42484 3000 42490 3052
rect 44726 3040 44732 3052
rect 44687 3012 44732 3040
rect 44726 3000 44732 3012
rect 44784 3000 44790 3052
rect 47857 3043 47915 3049
rect 47857 3009 47869 3043
rect 47903 3040 47915 3043
rect 49602 3040 49608 3052
rect 47903 3012 49608 3040
rect 47903 3009 47915 3012
rect 47857 3003 47915 3009
rect 49602 3000 49608 3012
rect 49660 3000 49666 3052
rect 8987 2944 12296 2972
rect 8987 2941 8999 2944
rect 8941 2935 8999 2941
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 12621 2975 12679 2981
rect 12492 2944 12537 2972
rect 12492 2932 12498 2944
rect 12621 2941 12633 2975
rect 12667 2972 12679 2975
rect 12710 2972 12716 2984
rect 12667 2944 12716 2972
rect 12667 2941 12679 2944
rect 12621 2935 12679 2941
rect 12710 2932 12716 2944
rect 12768 2932 12774 2984
rect 12894 2972 12900 2984
rect 12855 2944 12900 2972
rect 12894 2932 12900 2944
rect 12952 2932 12958 2984
rect 17586 2972 17592 2984
rect 13004 2944 17592 2972
rect 7098 2904 7104 2916
rect 6564 2876 7104 2904
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 10962 2864 10968 2916
rect 11020 2904 11026 2916
rect 13004 2904 13032 2944
rect 17586 2932 17592 2944
rect 17644 2932 17650 2984
rect 18046 2972 18052 2984
rect 18007 2944 18052 2972
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 23842 2972 23848 2984
rect 23803 2944 23848 2972
rect 23842 2932 23848 2944
rect 23900 2932 23906 2984
rect 24118 2932 24124 2984
rect 24176 2972 24182 2984
rect 24176 2944 26648 2972
rect 24176 2932 24182 2944
rect 11020 2876 13032 2904
rect 11020 2864 11026 2876
rect 20438 2864 20444 2916
rect 20496 2904 20502 2916
rect 26620 2904 26648 2944
rect 26694 2932 26700 2984
rect 26752 2972 26758 2984
rect 31202 2972 31208 2984
rect 26752 2944 31208 2972
rect 26752 2932 26758 2944
rect 31202 2932 31208 2944
rect 31260 2932 31266 2984
rect 31294 2932 31300 2984
rect 31352 2972 31358 2984
rect 33502 2972 33508 2984
rect 31352 2944 31397 2972
rect 33463 2944 33508 2972
rect 31352 2932 31358 2944
rect 33502 2932 33508 2944
rect 33560 2932 33566 2984
rect 34514 2932 34520 2984
rect 34572 2972 34578 2984
rect 38010 2972 38016 2984
rect 34572 2944 38016 2972
rect 34572 2932 34578 2944
rect 38010 2932 38016 2944
rect 38068 2932 38074 2984
rect 38746 2972 38752 2984
rect 38707 2944 38752 2972
rect 38746 2932 38752 2944
rect 38804 2932 38810 2984
rect 39942 2972 39948 2984
rect 39903 2944 39948 2972
rect 39942 2932 39948 2944
rect 40000 2932 40006 2984
rect 41601 2975 41659 2981
rect 41601 2941 41613 2975
rect 41647 2972 41659 2975
rect 42613 2975 42671 2981
rect 42613 2972 42625 2975
rect 41647 2944 42625 2972
rect 41647 2941 41659 2944
rect 41601 2935 41659 2941
rect 42613 2941 42625 2944
rect 42659 2941 42671 2975
rect 42613 2935 42671 2941
rect 42702 2932 42708 2984
rect 42760 2972 42766 2984
rect 42889 2975 42947 2981
rect 42889 2972 42901 2975
rect 42760 2944 42901 2972
rect 42760 2932 42766 2944
rect 42889 2941 42901 2944
rect 42935 2941 42947 2975
rect 42889 2935 42947 2941
rect 45094 2932 45100 2984
rect 45152 2972 45158 2984
rect 45189 2975 45247 2981
rect 45189 2972 45201 2975
rect 45152 2944 45201 2972
rect 45152 2932 45158 2944
rect 45189 2941 45201 2944
rect 45235 2941 45247 2975
rect 45189 2935 45247 2941
rect 32214 2904 32220 2916
rect 20496 2876 26556 2904
rect 26620 2876 32220 2904
rect 20496 2864 20502 2876
rect 2056 2808 5028 2836
rect 5810 2796 5816 2848
rect 5868 2836 5874 2848
rect 7006 2836 7012 2848
rect 5868 2808 7012 2836
rect 5868 2796 5874 2808
rect 7006 2796 7012 2808
rect 7064 2796 7070 2848
rect 11514 2796 11520 2848
rect 11572 2836 11578 2848
rect 18138 2836 18144 2848
rect 11572 2808 18144 2836
rect 11572 2796 11578 2808
rect 18138 2796 18144 2808
rect 18196 2796 18202 2848
rect 22738 2796 22744 2848
rect 22796 2836 22802 2848
rect 22833 2839 22891 2845
rect 22833 2836 22845 2839
rect 22796 2808 22845 2836
rect 22796 2796 22802 2808
rect 22833 2805 22845 2808
rect 22879 2805 22891 2839
rect 26142 2836 26148 2848
rect 26103 2808 26148 2836
rect 22833 2799 22891 2805
rect 26142 2796 26148 2808
rect 26200 2796 26206 2848
rect 26528 2836 26556 2876
rect 32214 2864 32220 2876
rect 32272 2864 32278 2916
rect 48041 2907 48099 2913
rect 48041 2904 48053 2907
rect 35866 2876 48053 2904
rect 35866 2836 35894 2876
rect 48041 2873 48053 2876
rect 48087 2873 48099 2907
rect 48041 2867 48099 2873
rect 26528 2808 35894 2836
rect 41874 2796 41880 2848
rect 41932 2836 41938 2848
rect 42702 2836 42708 2848
rect 41932 2808 42708 2836
rect 41932 2796 41938 2808
rect 42702 2796 42708 2808
rect 42760 2796 42766 2848
rect 1104 2746 48852 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 48852 2746
rect 1104 2672 48852 2694
rect 3970 2632 3976 2644
rect 3931 2604 3976 2632
rect 3970 2592 3976 2604
rect 4028 2592 4034 2644
rect 4062 2592 4068 2644
rect 4120 2632 4126 2644
rect 9122 2632 9128 2644
rect 4120 2604 9128 2632
rect 4120 2592 4126 2604
rect 9122 2592 9128 2604
rect 9180 2592 9186 2644
rect 12434 2592 12440 2644
rect 12492 2632 12498 2644
rect 12713 2635 12771 2641
rect 12713 2632 12725 2635
rect 12492 2604 12725 2632
rect 12492 2592 12498 2604
rect 12713 2601 12725 2604
rect 12759 2601 12771 2635
rect 12713 2595 12771 2601
rect 13170 2592 13176 2644
rect 13228 2632 13234 2644
rect 13357 2635 13415 2641
rect 13357 2632 13369 2635
rect 13228 2604 13369 2632
rect 13228 2592 13234 2604
rect 13357 2601 13369 2604
rect 13403 2601 13415 2635
rect 13357 2595 13415 2601
rect 21634 2592 21640 2644
rect 21692 2632 21698 2644
rect 46842 2632 46848 2644
rect 21692 2604 46848 2632
rect 21692 2592 21698 2604
rect 46842 2592 46848 2604
rect 46900 2592 46906 2644
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 7190 2564 7196 2576
rect 1360 2536 1900 2564
rect 1360 2524 1366 2536
rect 1397 2499 1455 2505
rect 1397 2465 1409 2499
rect 1443 2496 1455 2499
rect 1578 2496 1584 2508
rect 1443 2468 1584 2496
rect 1443 2465 1455 2468
rect 1397 2459 1455 2465
rect 1578 2456 1584 2468
rect 1636 2456 1642 2508
rect 1872 2505 1900 2536
rect 6380 2536 7196 2564
rect 6380 2505 6408 2536
rect 7190 2524 7196 2536
rect 7248 2524 7254 2576
rect 17773 2567 17831 2573
rect 17773 2533 17785 2567
rect 17819 2564 17831 2567
rect 20162 2564 20168 2576
rect 17819 2536 20168 2564
rect 17819 2533 17831 2536
rect 17773 2527 17831 2533
rect 20162 2524 20168 2536
rect 20220 2524 20226 2576
rect 20346 2564 20352 2576
rect 20307 2536 20352 2564
rect 20346 2524 20352 2536
rect 20404 2524 20410 2576
rect 21266 2524 21272 2576
rect 21324 2564 21330 2576
rect 21324 2536 22324 2564
rect 21324 2524 21330 2536
rect 1857 2499 1915 2505
rect 1857 2465 1869 2499
rect 1903 2465 1915 2499
rect 1857 2459 1915 2465
rect 6365 2499 6423 2505
rect 6365 2465 6377 2499
rect 6411 2465 6423 2499
rect 6365 2459 6423 2465
rect 6549 2499 6607 2505
rect 6549 2465 6561 2499
rect 6595 2496 6607 2499
rect 6914 2496 6920 2508
rect 6595 2468 6920 2496
rect 6595 2465 6607 2468
rect 6549 2459 6607 2465
rect 6914 2456 6920 2468
rect 6972 2456 6978 2508
rect 7006 2456 7012 2508
rect 7064 2496 7070 2508
rect 7064 2468 7109 2496
rect 7064 2456 7070 2468
rect 7466 2456 7472 2508
rect 7524 2496 7530 2508
rect 8941 2499 8999 2505
rect 8941 2496 8953 2499
rect 7524 2468 8953 2496
rect 7524 2456 7530 2468
rect 8941 2465 8953 2468
rect 8987 2465 8999 2499
rect 8941 2459 8999 2465
rect 9217 2499 9275 2505
rect 9217 2465 9229 2499
rect 9263 2496 9275 2499
rect 15194 2496 15200 2508
rect 9263 2468 15200 2496
rect 9263 2465 9275 2468
rect 9217 2459 9275 2465
rect 15194 2456 15200 2468
rect 15252 2456 15258 2508
rect 20990 2456 20996 2508
rect 21048 2496 21054 2508
rect 22296 2505 22324 2536
rect 24118 2524 24124 2576
rect 24176 2564 24182 2576
rect 25866 2564 25872 2576
rect 24176 2536 24992 2564
rect 25827 2536 25872 2564
rect 24176 2524 24182 2536
rect 21821 2499 21879 2505
rect 21821 2496 21833 2499
rect 21048 2468 21833 2496
rect 21048 2456 21054 2468
rect 21821 2465 21833 2468
rect 21867 2465 21879 2499
rect 21821 2459 21879 2465
rect 22281 2499 22339 2505
rect 22281 2465 22293 2499
rect 22327 2465 22339 2499
rect 22281 2459 22339 2465
rect 23934 2456 23940 2508
rect 23992 2496 23998 2508
rect 24857 2499 24915 2505
rect 24857 2496 24869 2499
rect 23992 2468 24869 2496
rect 23992 2456 23998 2468
rect 24857 2465 24869 2468
rect 24903 2465 24915 2499
rect 24964 2496 24992 2536
rect 25866 2524 25872 2536
rect 25924 2524 25930 2576
rect 27246 2564 27252 2576
rect 27207 2536 27252 2564
rect 27246 2524 27252 2536
rect 27304 2524 27310 2576
rect 30466 2564 30472 2576
rect 29748 2536 30472 2564
rect 29748 2505 29776 2536
rect 30466 2524 30472 2536
rect 30524 2524 30530 2576
rect 33134 2564 33140 2576
rect 33095 2536 33140 2564
rect 33134 2524 33140 2536
rect 33192 2524 33198 2576
rect 35066 2564 35072 2576
rect 35027 2536 35072 2564
rect 35066 2524 35072 2536
rect 35124 2524 35130 2576
rect 35342 2524 35348 2576
rect 35400 2564 35406 2576
rect 36173 2567 36231 2573
rect 36173 2564 36185 2567
rect 35400 2536 36185 2564
rect 35400 2524 35406 2536
rect 36173 2533 36185 2536
rect 36219 2533 36231 2567
rect 36173 2527 36231 2533
rect 38654 2524 38660 2576
rect 38712 2564 38718 2576
rect 38712 2536 38792 2564
rect 38712 2524 38718 2536
rect 28077 2499 28135 2505
rect 28077 2496 28089 2499
rect 24964 2468 28089 2496
rect 24857 2459 24915 2465
rect 28077 2465 28089 2468
rect 28123 2465 28135 2499
rect 28077 2459 28135 2465
rect 29733 2499 29791 2505
rect 29733 2465 29745 2499
rect 29779 2465 29791 2499
rect 29733 2459 29791 2465
rect 29917 2499 29975 2505
rect 29917 2465 29929 2499
rect 29963 2496 29975 2499
rect 30282 2496 30288 2508
rect 29963 2468 30288 2496
rect 29963 2465 29975 2468
rect 29917 2459 29975 2465
rect 30282 2456 30288 2468
rect 30340 2456 30346 2508
rect 30926 2496 30932 2508
rect 30887 2468 30932 2496
rect 30926 2456 30932 2468
rect 30984 2456 30990 2508
rect 38764 2505 38792 2536
rect 38749 2499 38807 2505
rect 38749 2465 38761 2499
rect 38795 2465 38807 2499
rect 38749 2459 38807 2465
rect 45189 2499 45247 2505
rect 45189 2465 45201 2499
rect 45235 2496 45247 2499
rect 45830 2496 45836 2508
rect 45235 2468 45836 2496
rect 45235 2465 45247 2468
rect 45189 2459 45247 2465
rect 45830 2456 45836 2468
rect 45888 2456 45894 2508
rect 4522 2388 4528 2440
rect 4580 2428 4586 2440
rect 4617 2431 4675 2437
rect 4617 2428 4629 2431
rect 4580 2400 4629 2428
rect 4580 2388 4586 2400
rect 4617 2397 4629 2400
rect 4663 2397 4675 2431
rect 4617 2391 4675 2397
rect 14737 2431 14795 2437
rect 14737 2397 14749 2431
rect 14783 2428 14795 2431
rect 20530 2428 20536 2440
rect 14783 2400 20536 2428
rect 14783 2397 14795 2400
rect 14737 2391 14795 2397
rect 20530 2388 20536 2400
rect 20588 2388 20594 2440
rect 24486 2388 24492 2440
rect 24544 2428 24550 2440
rect 24581 2431 24639 2437
rect 24581 2428 24593 2431
rect 24544 2400 24593 2428
rect 24544 2388 24550 2400
rect 24581 2397 24593 2400
rect 24627 2397 24639 2431
rect 24581 2391 24639 2397
rect 25130 2388 25136 2440
rect 25188 2428 25194 2440
rect 26053 2431 26111 2437
rect 26053 2428 26065 2431
rect 25188 2400 26065 2428
rect 25188 2388 25194 2400
rect 26053 2397 26065 2400
rect 26099 2397 26111 2431
rect 27062 2428 27068 2440
rect 27023 2400 27068 2428
rect 26053 2391 26111 2397
rect 27062 2388 27068 2400
rect 27120 2388 27126 2440
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27764 2400 27813 2428
rect 27764 2388 27770 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 32858 2388 32864 2440
rect 32916 2428 32922 2440
rect 32953 2431 33011 2437
rect 32953 2428 32965 2431
rect 32916 2400 32965 2428
rect 32916 2388 32922 2400
rect 32953 2397 32965 2400
rect 32999 2397 33011 2431
rect 32953 2391 33011 2397
rect 33060 2400 34284 2428
rect 1581 2363 1639 2369
rect 1581 2329 1593 2363
rect 1627 2360 1639 2363
rect 2866 2360 2872 2372
rect 1627 2332 2872 2360
rect 1627 2329 1639 2332
rect 1581 2323 1639 2329
rect 2866 2320 2872 2332
rect 2924 2320 2930 2372
rect 8386 2320 8392 2372
rect 8444 2360 8450 2372
rect 10321 2363 10379 2369
rect 10321 2360 10333 2363
rect 8444 2332 10333 2360
rect 8444 2320 8450 2332
rect 10321 2329 10333 2332
rect 10367 2329 10379 2363
rect 10321 2323 10379 2329
rect 14182 2320 14188 2372
rect 14240 2360 14246 2372
rect 14553 2363 14611 2369
rect 14553 2360 14565 2363
rect 14240 2332 14565 2360
rect 14240 2320 14246 2332
rect 14553 2329 14565 2332
rect 14599 2329 14611 2363
rect 14553 2323 14611 2329
rect 17402 2320 17408 2372
rect 17460 2360 17466 2372
rect 17589 2363 17647 2369
rect 17589 2360 17601 2363
rect 17460 2332 17601 2360
rect 17460 2320 17466 2332
rect 17589 2329 17601 2332
rect 17635 2329 17647 2363
rect 17589 2323 17647 2329
rect 19978 2320 19984 2372
rect 20036 2360 20042 2372
rect 20165 2363 20223 2369
rect 20165 2360 20177 2363
rect 20036 2332 20177 2360
rect 20036 2320 20042 2332
rect 20165 2329 20177 2332
rect 20211 2329 20223 2363
rect 20165 2323 20223 2329
rect 21082 2320 21088 2372
rect 21140 2360 21146 2372
rect 22005 2363 22063 2369
rect 22005 2360 22017 2363
rect 21140 2332 22017 2360
rect 21140 2320 21146 2332
rect 22005 2329 22017 2332
rect 22051 2329 22063 2363
rect 22005 2323 22063 2329
rect 25774 2320 25780 2372
rect 25832 2360 25838 2372
rect 33060 2360 33088 2400
rect 25832 2332 33088 2360
rect 33965 2363 34023 2369
rect 25832 2320 25838 2332
rect 33965 2329 33977 2363
rect 34011 2360 34023 2363
rect 34146 2360 34152 2372
rect 34011 2332 34152 2360
rect 34011 2329 34023 2332
rect 33965 2323 34023 2329
rect 34146 2320 34152 2332
rect 34204 2320 34210 2372
rect 4798 2292 4804 2304
rect 4759 2264 4804 2292
rect 4798 2252 4804 2264
rect 4856 2252 4862 2304
rect 10594 2292 10600 2304
rect 10555 2264 10600 2292
rect 10594 2252 10600 2264
rect 10652 2252 10658 2304
rect 23014 2252 23020 2304
rect 23072 2292 23078 2304
rect 34057 2295 34115 2301
rect 34057 2292 34069 2295
rect 23072 2264 34069 2292
rect 23072 2252 23078 2264
rect 34057 2261 34069 2264
rect 34103 2261 34115 2295
rect 34256 2292 34284 2400
rect 34790 2388 34796 2440
rect 34848 2428 34854 2440
rect 34885 2431 34943 2437
rect 34885 2428 34897 2431
rect 34848 2400 34897 2428
rect 34848 2388 34854 2400
rect 34885 2397 34897 2400
rect 34931 2397 34943 2431
rect 34885 2391 34943 2397
rect 36078 2388 36084 2440
rect 36136 2428 36142 2440
rect 36357 2431 36415 2437
rect 36357 2428 36369 2431
rect 36136 2400 36369 2428
rect 36136 2388 36142 2400
rect 36357 2397 36369 2400
rect 36403 2397 36415 2431
rect 36357 2391 36415 2397
rect 38473 2431 38531 2437
rect 38473 2397 38485 2431
rect 38519 2428 38531 2431
rect 38654 2428 38660 2440
rect 38519 2400 38660 2428
rect 38519 2397 38531 2400
rect 38473 2391 38531 2397
rect 38654 2388 38660 2400
rect 38712 2388 38718 2440
rect 44453 2431 44511 2437
rect 44453 2428 44465 2431
rect 38764 2400 44465 2428
rect 38102 2320 38108 2372
rect 38160 2360 38166 2372
rect 38764 2360 38792 2400
rect 44453 2397 44465 2400
rect 44499 2397 44511 2431
rect 44453 2391 44511 2397
rect 47029 2431 47087 2437
rect 47029 2397 47041 2431
rect 47075 2428 47087 2431
rect 48314 2428 48320 2440
rect 47075 2400 48320 2428
rect 47075 2397 47087 2400
rect 47029 2391 47087 2397
rect 48314 2388 48320 2400
rect 48372 2388 48378 2440
rect 38160 2332 38792 2360
rect 38160 2320 38166 2332
rect 43162 2320 43168 2372
rect 43220 2360 43226 2372
rect 43349 2363 43407 2369
rect 43349 2360 43361 2363
rect 43220 2332 43361 2360
rect 43220 2320 43226 2332
rect 43349 2329 43361 2332
rect 43395 2329 43407 2363
rect 43349 2323 43407 2329
rect 44269 2363 44327 2369
rect 44269 2329 44281 2363
rect 44315 2360 44327 2363
rect 45373 2363 45431 2369
rect 44315 2332 44956 2360
rect 44315 2329 44327 2332
rect 44269 2323 44327 2329
rect 43441 2295 43499 2301
rect 43441 2292 43453 2295
rect 34256 2264 43453 2292
rect 34057 2255 34115 2261
rect 43441 2261 43453 2264
rect 43487 2261 43499 2295
rect 44928 2292 44956 2332
rect 45373 2329 45385 2363
rect 45419 2360 45431 2363
rect 46934 2360 46940 2372
rect 45419 2332 46940 2360
rect 45419 2329 45431 2332
rect 45373 2323 45431 2329
rect 46934 2320 46940 2332
rect 46992 2320 46998 2372
rect 47762 2360 47768 2372
rect 47723 2332 47768 2360
rect 47762 2320 47768 2332
rect 47820 2320 47826 2372
rect 45738 2292 45744 2304
rect 44928 2264 45744 2292
rect 43441 2255 43499 2261
rect 45738 2252 45744 2264
rect 45796 2252 45802 2304
rect 47854 2292 47860 2304
rect 47815 2264 47860 2292
rect 47854 2252 47860 2264
rect 47912 2252 47918 2304
rect 1104 2202 48852 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 48852 2202
rect 1104 2128 48852 2150
rect 21818 2048 21824 2100
rect 21876 2088 21882 2100
rect 27246 2088 27252 2100
rect 21876 2060 27252 2088
rect 21876 2048 21882 2060
rect 27246 2048 27252 2060
rect 27304 2048 27310 2100
rect 21174 1980 21180 2032
rect 21232 2020 21238 2032
rect 33134 2020 33140 2032
rect 21232 1992 33140 2020
rect 21232 1980 21238 1992
rect 33134 1980 33140 1992
rect 33192 1980 33198 2032
rect 10594 1912 10600 1964
rect 10652 1952 10658 1964
rect 28718 1952 28724 1964
rect 10652 1924 28724 1952
rect 10652 1912 10658 1924
rect 28718 1912 28724 1924
rect 28776 1912 28782 1964
rect 26510 1844 26516 1896
rect 26568 1884 26574 1896
rect 47854 1884 47860 1896
rect 26568 1856 47860 1884
rect 26568 1844 26574 1856
rect 47854 1844 47860 1856
rect 47912 1844 47918 1896
rect 12250 1232 12256 1284
rect 12308 1272 12314 1284
rect 12802 1272 12808 1284
rect 12308 1244 12808 1272
rect 12308 1232 12314 1244
rect 12802 1232 12808 1244
rect 12860 1232 12866 1284
<< via1 >>
rect 4068 49716 4120 49768
rect 5632 49716 5684 49768
rect 37004 49716 37056 49768
rect 45560 49716 45612 49768
rect 4214 49478 4266 49530
rect 4278 49478 4330 49530
rect 4342 49478 4394 49530
rect 4406 49478 4458 49530
rect 4470 49478 4522 49530
rect 34934 49478 34986 49530
rect 34998 49478 35050 49530
rect 35062 49478 35114 49530
rect 35126 49478 35178 49530
rect 35190 49478 35242 49530
rect 6920 49240 6972 49292
rect 7104 49283 7156 49292
rect 7104 49249 7113 49283
rect 7113 49249 7147 49283
rect 7147 49249 7156 49283
rect 7104 49240 7156 49249
rect 7748 49240 7800 49292
rect 12716 49283 12768 49292
rect 12716 49249 12725 49283
rect 12725 49249 12759 49283
rect 12759 49249 12768 49283
rect 12716 49240 12768 49249
rect 14464 49240 14516 49292
rect 664 49172 716 49224
rect 3608 49172 3660 49224
rect 4620 49172 4672 49224
rect 8944 49215 8996 49224
rect 8944 49181 8953 49215
rect 8953 49181 8987 49215
rect 8987 49181 8996 49215
rect 8944 49172 8996 49181
rect 11612 49172 11664 49224
rect 2780 49147 2832 49156
rect 2780 49113 2789 49147
rect 2789 49113 2823 49147
rect 2823 49113 2832 49147
rect 2780 49104 2832 49113
rect 2964 49147 3016 49156
rect 2964 49113 2973 49147
rect 2973 49113 3007 49147
rect 3007 49113 3016 49147
rect 2964 49104 3016 49113
rect 7380 49104 7432 49156
rect 8484 49104 8536 49156
rect 13820 49172 13872 49224
rect 16580 49240 16632 49292
rect 24124 49308 24176 49360
rect 29920 49308 29972 49360
rect 33508 49308 33560 49360
rect 34428 49308 34480 49360
rect 22560 49283 22612 49292
rect 22560 49249 22569 49283
rect 22569 49249 22603 49283
rect 22603 49249 22612 49283
rect 22560 49240 22612 49249
rect 30472 49240 30524 49292
rect 30932 49283 30984 49292
rect 30932 49249 30941 49283
rect 30941 49249 30975 49283
rect 30975 49249 30984 49283
rect 30932 49240 30984 49249
rect 43168 49283 43220 49292
rect 43168 49249 43177 49283
rect 43177 49249 43211 49283
rect 43211 49249 43220 49283
rect 43168 49240 43220 49249
rect 45192 49240 45244 49292
rect 17960 49172 18012 49224
rect 19432 49215 19484 49224
rect 19432 49181 19441 49215
rect 19441 49181 19475 49215
rect 19475 49181 19484 49215
rect 19432 49172 19484 49181
rect 20076 49215 20128 49224
rect 20076 49181 20085 49215
rect 20085 49181 20119 49215
rect 20119 49181 20128 49215
rect 20076 49172 20128 49181
rect 21640 49172 21692 49224
rect 21824 49215 21876 49224
rect 21824 49181 21833 49215
rect 21833 49181 21867 49215
rect 21867 49181 21876 49215
rect 21824 49172 21876 49181
rect 23848 49172 23900 49224
rect 25964 49215 26016 49224
rect 25964 49181 25973 49215
rect 25973 49181 26007 49215
rect 26007 49181 26016 49215
rect 25964 49172 26016 49181
rect 26424 49172 26476 49224
rect 27988 49172 28040 49224
rect 29000 49172 29052 49224
rect 31944 49172 31996 49224
rect 33508 49172 33560 49224
rect 34888 49172 34940 49224
rect 36176 49215 36228 49224
rect 36176 49181 36185 49215
rect 36185 49181 36219 49215
rect 36219 49181 36228 49215
rect 36176 49172 36228 49181
rect 38200 49215 38252 49224
rect 38200 49181 38209 49215
rect 38209 49181 38243 49215
rect 38243 49181 38252 49215
rect 38200 49172 38252 49181
rect 43996 49172 44048 49224
rect 47768 49215 47820 49224
rect 47768 49181 47777 49215
rect 47777 49181 47811 49215
rect 47811 49181 47820 49215
rect 47768 49172 47820 49181
rect 17224 49104 17276 49156
rect 20536 49104 20588 49156
rect 22284 49104 22336 49156
rect 27712 49104 27764 49156
rect 30656 49104 30708 49156
rect 40776 49147 40828 49156
rect 40776 49113 40785 49147
rect 40785 49113 40819 49147
rect 40819 49113 40828 49147
rect 40776 49104 40828 49113
rect 41696 49104 41748 49156
rect 41788 49104 41840 49156
rect 44088 49104 44140 49156
rect 1492 49036 1544 49088
rect 4620 49036 4672 49088
rect 5264 49079 5316 49088
rect 5264 49045 5273 49079
rect 5273 49045 5307 49079
rect 5307 49045 5316 49079
rect 5264 49036 5316 49045
rect 12072 49079 12124 49088
rect 12072 49045 12081 49079
rect 12081 49045 12115 49079
rect 12115 49045 12124 49079
rect 12072 49036 12124 49045
rect 14648 49079 14700 49088
rect 14648 49045 14657 49079
rect 14657 49045 14691 49079
rect 14691 49045 14700 49079
rect 14648 49036 14700 49045
rect 17592 49036 17644 49088
rect 20352 49036 20404 49088
rect 21088 49079 21140 49088
rect 21088 49045 21097 49079
rect 21097 49045 21131 49079
rect 21131 49045 21140 49079
rect 21088 49036 21140 49045
rect 22376 49036 22428 49088
rect 25412 49036 25464 49088
rect 32128 49036 32180 49088
rect 38016 49036 38068 49088
rect 40868 49079 40920 49088
rect 40868 49045 40877 49079
rect 40877 49045 40911 49079
rect 40911 49045 40920 49079
rect 40868 49036 40920 49045
rect 41604 49079 41656 49088
rect 41604 49045 41613 49079
rect 41613 49045 41647 49079
rect 41647 49045 41656 49079
rect 41604 49036 41656 49045
rect 47308 49036 47360 49088
rect 19574 48934 19626 48986
rect 19638 48934 19690 48986
rect 19702 48934 19754 48986
rect 19766 48934 19818 48986
rect 19830 48934 19882 48986
rect 41788 48875 41840 48884
rect 41788 48841 41797 48875
rect 41797 48841 41831 48875
rect 41831 48841 41840 48875
rect 41788 48832 41840 48841
rect 2872 48764 2924 48816
rect 5540 48764 5592 48816
rect 3056 48628 3108 48680
rect 4896 48628 4948 48680
rect 5632 48671 5684 48680
rect 5632 48637 5641 48671
rect 5641 48637 5675 48671
rect 5675 48637 5684 48671
rect 5632 48628 5684 48637
rect 6368 48671 6420 48680
rect 6368 48637 6377 48671
rect 6377 48637 6411 48671
rect 6411 48637 6420 48671
rect 6368 48628 6420 48637
rect 7564 48628 7616 48680
rect 10508 48764 10560 48816
rect 34796 48764 34848 48816
rect 36728 48807 36780 48816
rect 36728 48773 36737 48807
rect 36737 48773 36771 48807
rect 36771 48773 36780 48807
rect 36728 48764 36780 48773
rect 48320 48832 48372 48884
rect 47768 48807 47820 48816
rect 47768 48773 47777 48807
rect 47777 48773 47811 48807
rect 47811 48773 47820 48807
rect 47768 48764 47820 48773
rect 18052 48696 18104 48748
rect 21824 48696 21876 48748
rect 32128 48739 32180 48748
rect 32128 48705 32137 48739
rect 32137 48705 32171 48739
rect 32171 48705 32180 48739
rect 32128 48696 32180 48705
rect 34888 48739 34940 48748
rect 34888 48705 34897 48739
rect 34897 48705 34931 48739
rect 34931 48705 34940 48739
rect 34888 48696 34940 48705
rect 41696 48739 41748 48748
rect 41696 48705 41705 48739
rect 41705 48705 41739 48739
rect 41739 48705 41748 48739
rect 41696 48696 41748 48705
rect 9128 48671 9180 48680
rect 9128 48637 9137 48671
rect 9137 48637 9171 48671
rect 9171 48637 9180 48671
rect 9128 48628 9180 48637
rect 9680 48671 9732 48680
rect 9680 48637 9689 48671
rect 9689 48637 9723 48671
rect 9723 48637 9732 48671
rect 9680 48628 9732 48637
rect 12440 48671 12492 48680
rect 12440 48637 12449 48671
rect 12449 48637 12483 48671
rect 12483 48637 12492 48671
rect 12440 48628 12492 48637
rect 12808 48628 12860 48680
rect 16856 48671 16908 48680
rect 4712 48560 4764 48612
rect 12532 48560 12584 48612
rect 16856 48637 16865 48671
rect 16865 48637 16899 48671
rect 16899 48637 16908 48671
rect 16856 48628 16908 48637
rect 17040 48628 17092 48680
rect 22652 48671 22704 48680
rect 22652 48637 22661 48671
rect 22661 48637 22695 48671
rect 22695 48637 22704 48671
rect 22652 48628 22704 48637
rect 23480 48671 23532 48680
rect 23480 48637 23489 48671
rect 23489 48637 23523 48671
rect 23523 48637 23532 48671
rect 23480 48628 23532 48637
rect 27252 48671 27304 48680
rect 27252 48637 27261 48671
rect 27261 48637 27295 48671
rect 27295 48637 27304 48671
rect 27252 48628 27304 48637
rect 27804 48671 27856 48680
rect 27804 48637 27813 48671
rect 27813 48637 27847 48671
rect 27847 48637 27856 48671
rect 27804 48628 27856 48637
rect 29276 48628 29328 48680
rect 29552 48671 29604 48680
rect 29552 48637 29561 48671
rect 29561 48637 29595 48671
rect 29595 48637 29604 48671
rect 29552 48628 29604 48637
rect 29828 48671 29880 48680
rect 29828 48637 29837 48671
rect 29837 48637 29871 48671
rect 29871 48637 29880 48671
rect 29828 48628 29880 48637
rect 32312 48671 32364 48680
rect 32312 48637 32321 48671
rect 32321 48637 32355 48671
rect 32355 48637 32364 48671
rect 32312 48628 32364 48637
rect 33140 48671 33192 48680
rect 33140 48637 33149 48671
rect 33149 48637 33183 48671
rect 33183 48637 33192 48671
rect 33140 48628 33192 48637
rect 39396 48671 39448 48680
rect 39396 48637 39405 48671
rect 39405 48637 39439 48671
rect 39439 48637 39448 48671
rect 39396 48628 39448 48637
rect 40040 48671 40092 48680
rect 40040 48637 40049 48671
rect 40049 48637 40083 48671
rect 40083 48637 40092 48671
rect 40040 48628 40092 48637
rect 41420 48628 41472 48680
rect 43076 48671 43128 48680
rect 43076 48637 43085 48671
rect 43085 48637 43119 48671
rect 43119 48637 43128 48671
rect 43076 48628 43128 48637
rect 44824 48628 44876 48680
rect 45376 48671 45428 48680
rect 45376 48637 45385 48671
rect 45385 48637 45419 48671
rect 45419 48637 45428 48671
rect 45376 48628 45428 48637
rect 45744 48671 45796 48680
rect 45744 48637 45753 48671
rect 45753 48637 45787 48671
rect 45787 48637 45796 48671
rect 45744 48628 45796 48637
rect 5356 48492 5408 48544
rect 11704 48535 11756 48544
rect 11704 48501 11713 48535
rect 11713 48501 11747 48535
rect 11747 48501 11756 48535
rect 11704 48492 11756 48501
rect 14924 48535 14976 48544
rect 14924 48501 14933 48535
rect 14933 48501 14967 48535
rect 14967 48501 14976 48535
rect 14924 48492 14976 48501
rect 18052 48492 18104 48544
rect 20444 48535 20496 48544
rect 20444 48501 20453 48535
rect 20453 48501 20487 48535
rect 20487 48501 20496 48535
rect 20444 48492 20496 48501
rect 24952 48535 25004 48544
rect 24952 48501 24961 48535
rect 24961 48501 24995 48535
rect 24995 48501 25004 48535
rect 24952 48492 25004 48501
rect 26700 48492 26752 48544
rect 47124 48492 47176 48544
rect 4214 48390 4266 48442
rect 4278 48390 4330 48442
rect 4342 48390 4394 48442
rect 4406 48390 4458 48442
rect 4470 48390 4522 48442
rect 34934 48390 34986 48442
rect 34998 48390 35050 48442
rect 35062 48390 35114 48442
rect 35126 48390 35178 48442
rect 35190 48390 35242 48442
rect 3424 48288 3476 48340
rect 6644 48288 6696 48340
rect 12440 48288 12492 48340
rect 12808 48288 12860 48340
rect 22652 48288 22704 48340
rect 20 48220 72 48272
rect 2780 48220 2832 48272
rect 3976 48220 4028 48272
rect 7380 48263 7432 48272
rect 1308 48152 1360 48204
rect 5540 48152 5592 48204
rect 7380 48229 7389 48263
rect 7389 48229 7423 48263
rect 7423 48229 7432 48263
rect 7380 48220 7432 48229
rect 7564 48220 7616 48272
rect 17408 48220 17460 48272
rect 9128 48152 9180 48204
rect 11704 48152 11756 48204
rect 14924 48152 14976 48204
rect 15016 48152 15068 48204
rect 17960 48152 18012 48204
rect 20444 48152 20496 48204
rect 20628 48152 20680 48204
rect 3792 48127 3844 48136
rect 3792 48093 3801 48127
rect 3801 48093 3835 48127
rect 3835 48093 3844 48127
rect 3792 48084 3844 48093
rect 7196 48084 7248 48136
rect 7932 48127 7984 48136
rect 7932 48093 7941 48127
rect 7941 48093 7975 48127
rect 7975 48093 7984 48127
rect 7932 48084 7984 48093
rect 24492 48220 24544 48272
rect 29552 48288 29604 48340
rect 34796 48331 34848 48340
rect 34796 48297 34805 48331
rect 34805 48297 34839 48331
rect 34839 48297 34848 48331
rect 34796 48288 34848 48297
rect 39396 48288 39448 48340
rect 30656 48263 30708 48272
rect 24952 48152 25004 48204
rect 26700 48195 26752 48204
rect 26700 48161 26709 48195
rect 26709 48161 26743 48195
rect 26743 48161 26752 48195
rect 26700 48152 26752 48161
rect 27068 48152 27120 48204
rect 23664 48127 23716 48136
rect 1584 48059 1636 48068
rect 1584 48025 1593 48059
rect 1593 48025 1627 48059
rect 1627 48025 1636 48059
rect 1584 48016 1636 48025
rect 4988 48016 5040 48068
rect 10048 48059 10100 48068
rect 10048 48025 10057 48059
rect 10057 48025 10091 48059
rect 10091 48025 10100 48059
rect 10048 48016 10100 48025
rect 10324 48016 10376 48068
rect 3884 47948 3936 48000
rect 4068 47948 4120 48000
rect 23664 48093 23673 48127
rect 23673 48093 23707 48127
rect 23707 48093 23716 48127
rect 23664 48084 23716 48093
rect 29552 48127 29604 48136
rect 29552 48093 29561 48127
rect 29561 48093 29595 48127
rect 29595 48093 29604 48127
rect 29552 48084 29604 48093
rect 30656 48229 30665 48263
rect 30665 48229 30699 48263
rect 30699 48229 30708 48263
rect 30656 48220 30708 48229
rect 36636 48220 36688 48272
rect 47032 48220 47084 48272
rect 49608 48220 49660 48272
rect 31944 48152 31996 48204
rect 32220 48195 32272 48204
rect 32220 48161 32229 48195
rect 32229 48161 32263 48195
rect 32263 48161 32272 48195
rect 32220 48152 32272 48161
rect 36176 48152 36228 48204
rect 36268 48195 36320 48204
rect 36268 48161 36277 48195
rect 36277 48161 36311 48195
rect 36311 48161 36320 48195
rect 42524 48195 42576 48204
rect 36268 48152 36320 48161
rect 42524 48161 42533 48195
rect 42533 48161 42567 48195
rect 42567 48161 42576 48195
rect 42524 48152 42576 48161
rect 46664 48152 46716 48204
rect 46848 48195 46900 48204
rect 46848 48161 46857 48195
rect 46857 48161 46891 48195
rect 46891 48161 46900 48195
rect 46848 48152 46900 48161
rect 30564 48127 30616 48136
rect 30564 48093 30573 48127
rect 30573 48093 30607 48127
rect 30607 48093 30616 48127
rect 30564 48084 30616 48093
rect 14372 48016 14424 48068
rect 17408 48016 17460 48068
rect 20260 48016 20312 48068
rect 16672 47948 16724 48000
rect 17132 47948 17184 48000
rect 23572 48016 23624 48068
rect 26332 48016 26384 48068
rect 31116 48016 31168 48068
rect 24032 47948 24084 48000
rect 33324 48084 33376 48136
rect 34612 48084 34664 48136
rect 43904 48127 43956 48136
rect 35900 48016 35952 48068
rect 33692 47991 33744 48000
rect 33692 47957 33701 47991
rect 33701 47957 33735 47991
rect 33735 47957 33744 47991
rect 33692 47948 33744 47957
rect 43904 48093 43913 48127
rect 43913 48093 43947 48127
rect 43947 48093 43956 48127
rect 43904 48084 43956 48093
rect 44456 48084 44508 48136
rect 41788 48016 41840 48068
rect 46480 48059 46532 48068
rect 46480 48025 46489 48059
rect 46489 48025 46523 48059
rect 46523 48025 46532 48059
rect 46480 48016 46532 48025
rect 44364 47948 44416 48000
rect 44916 47948 44968 48000
rect 19574 47846 19626 47898
rect 19638 47846 19690 47898
rect 19702 47846 19754 47898
rect 19766 47846 19818 47898
rect 19830 47846 19882 47898
rect 1584 47744 1636 47796
rect 4988 47787 5040 47796
rect 4988 47753 4997 47787
rect 4997 47753 5031 47787
rect 5031 47753 5040 47787
rect 4988 47744 5040 47753
rect 10048 47744 10100 47796
rect 10508 47787 10560 47796
rect 10508 47753 10517 47787
rect 10517 47753 10551 47787
rect 10551 47753 10560 47787
rect 10508 47744 10560 47753
rect 14372 47787 14424 47796
rect 14372 47753 14381 47787
rect 14381 47753 14415 47787
rect 14415 47753 14424 47787
rect 14372 47744 14424 47753
rect 16856 47744 16908 47796
rect 17408 47787 17460 47796
rect 17408 47753 17417 47787
rect 17417 47753 17451 47787
rect 17451 47753 17460 47787
rect 17408 47744 17460 47753
rect 20260 47787 20312 47796
rect 20260 47753 20269 47787
rect 20269 47753 20303 47787
rect 20303 47753 20312 47787
rect 20260 47744 20312 47753
rect 22284 47787 22336 47796
rect 22284 47753 22293 47787
rect 22293 47753 22327 47787
rect 22327 47753 22336 47787
rect 22284 47744 22336 47753
rect 26332 47787 26384 47796
rect 26332 47753 26341 47787
rect 26341 47753 26375 47787
rect 26375 47753 26384 47787
rect 26332 47744 26384 47753
rect 27252 47744 27304 47796
rect 31116 47787 31168 47796
rect 31116 47753 31125 47787
rect 31125 47753 31159 47787
rect 31159 47753 31168 47787
rect 31116 47744 31168 47753
rect 32312 47744 32364 47796
rect 6184 47676 6236 47728
rect 4804 47608 4856 47660
rect 6092 47608 6144 47660
rect 8944 47608 8996 47660
rect 14280 47651 14332 47660
rect 14280 47617 14289 47651
rect 14289 47617 14323 47651
rect 14323 47617 14332 47651
rect 14280 47608 14332 47617
rect 16672 47651 16724 47660
rect 16672 47617 16681 47651
rect 16681 47617 16715 47651
rect 16715 47617 16724 47651
rect 16672 47608 16724 47617
rect 17776 47608 17828 47660
rect 20168 47651 20220 47660
rect 20168 47617 20177 47651
rect 20177 47617 20211 47651
rect 20211 47617 20220 47651
rect 20168 47608 20220 47617
rect 23572 47676 23624 47728
rect 20996 47608 21048 47660
rect 22560 47608 22612 47660
rect 26516 47676 26568 47728
rect 41696 47744 41748 47796
rect 43076 47744 43128 47796
rect 33692 47719 33744 47728
rect 33692 47685 33701 47719
rect 33701 47685 33735 47719
rect 33735 47685 33744 47719
rect 33692 47676 33744 47685
rect 35900 47719 35952 47728
rect 35900 47685 35909 47719
rect 35909 47685 35943 47719
rect 35943 47685 35952 47719
rect 35900 47676 35952 47685
rect 27160 47608 27212 47660
rect 27988 47651 28040 47660
rect 27988 47617 27997 47651
rect 27997 47617 28031 47651
rect 28031 47617 28040 47651
rect 27988 47608 28040 47617
rect 30472 47651 30524 47660
rect 30472 47617 30481 47651
rect 30481 47617 30515 47651
rect 30515 47617 30524 47651
rect 30472 47608 30524 47617
rect 31024 47651 31076 47660
rect 31024 47617 31033 47651
rect 31033 47617 31067 47651
rect 31067 47617 31076 47651
rect 31024 47608 31076 47617
rect 32404 47651 32456 47660
rect 32404 47617 32413 47651
rect 32413 47617 32447 47651
rect 32447 47617 32456 47651
rect 32404 47608 32456 47617
rect 33508 47651 33560 47660
rect 33508 47617 33517 47651
rect 33517 47617 33551 47651
rect 33551 47617 33560 47651
rect 33508 47608 33560 47617
rect 35808 47651 35860 47660
rect 35808 47617 35817 47651
rect 35817 47617 35851 47651
rect 35851 47617 35860 47651
rect 35808 47608 35860 47617
rect 41420 47608 41472 47660
rect 45560 47676 45612 47728
rect 47768 47719 47820 47728
rect 47768 47685 47777 47719
rect 47777 47685 47811 47719
rect 47811 47685 47820 47719
rect 47768 47676 47820 47685
rect 1952 47583 2004 47592
rect 1952 47549 1961 47583
rect 1961 47549 1995 47583
rect 1995 47549 2004 47583
rect 1952 47540 2004 47549
rect 2872 47540 2924 47592
rect 3148 47583 3200 47592
rect 3148 47549 3157 47583
rect 3157 47549 3191 47583
rect 3191 47549 3200 47583
rect 3148 47540 3200 47549
rect 6552 47583 6604 47592
rect 6552 47549 6561 47583
rect 6561 47549 6595 47583
rect 6595 47549 6604 47583
rect 6552 47540 6604 47549
rect 6644 47540 6696 47592
rect 26424 47540 26476 47592
rect 28172 47583 28224 47592
rect 28172 47549 28181 47583
rect 28181 47549 28215 47583
rect 28215 47549 28224 47583
rect 28172 47540 28224 47549
rect 28448 47583 28500 47592
rect 28448 47549 28457 47583
rect 28457 47549 28491 47583
rect 28491 47549 28500 47583
rect 28448 47540 28500 47549
rect 34704 47583 34756 47592
rect 34704 47549 34713 47583
rect 34713 47549 34747 47583
rect 34747 47549 34756 47583
rect 34704 47540 34756 47549
rect 42708 47608 42760 47660
rect 42800 47540 42852 47592
rect 45100 47583 45152 47592
rect 17408 47472 17460 47524
rect 34612 47472 34664 47524
rect 6644 47404 6696 47456
rect 20536 47404 20588 47456
rect 20996 47404 21048 47456
rect 31024 47404 31076 47456
rect 31300 47404 31352 47456
rect 45100 47549 45109 47583
rect 45109 47549 45143 47583
rect 45143 47549 45152 47583
rect 45100 47540 45152 47549
rect 45284 47583 45336 47592
rect 45284 47549 45293 47583
rect 45293 47549 45327 47583
rect 45327 47549 45336 47583
rect 45284 47540 45336 47549
rect 46572 47583 46624 47592
rect 46572 47549 46581 47583
rect 46581 47549 46615 47583
rect 46615 47549 46624 47583
rect 46572 47540 46624 47549
rect 46572 47404 46624 47456
rect 47584 47404 47636 47456
rect 4214 47302 4266 47354
rect 4278 47302 4330 47354
rect 4342 47302 4394 47354
rect 4406 47302 4458 47354
rect 4470 47302 4522 47354
rect 34934 47302 34986 47354
rect 34998 47302 35050 47354
rect 35062 47302 35114 47354
rect 35126 47302 35178 47354
rect 35190 47302 35242 47354
rect 3056 47200 3108 47252
rect 4896 47200 4948 47252
rect 5540 47243 5592 47252
rect 5540 47209 5549 47243
rect 5549 47209 5583 47243
rect 5583 47209 5592 47243
rect 5540 47200 5592 47209
rect 6552 47200 6604 47252
rect 6920 47200 6972 47252
rect 8484 47200 8536 47252
rect 10968 47200 11020 47252
rect 13268 47200 13320 47252
rect 14280 47200 14332 47252
rect 24032 47200 24084 47252
rect 28172 47200 28224 47252
rect 3608 47132 3660 47184
rect 1860 47107 1912 47116
rect 1860 47073 1869 47107
rect 1869 47073 1903 47107
rect 1903 47073 1912 47107
rect 1860 47064 1912 47073
rect 17132 47132 17184 47184
rect 3332 46996 3384 47048
rect 6092 46996 6144 47048
rect 7748 47039 7800 47048
rect 1584 46971 1636 46980
rect 1584 46937 1593 46971
rect 1593 46937 1627 46971
rect 1627 46937 1636 46971
rect 1584 46928 1636 46937
rect 7748 47005 7757 47039
rect 7757 47005 7791 47039
rect 7791 47005 7800 47039
rect 7748 46996 7800 47005
rect 7932 46996 7984 47048
rect 20536 47107 20588 47116
rect 20536 47073 20545 47107
rect 20545 47073 20579 47107
rect 20579 47073 20588 47107
rect 20536 47064 20588 47073
rect 29552 47132 29604 47184
rect 42340 47200 42392 47252
rect 45284 47200 45336 47252
rect 35808 47132 35860 47184
rect 20352 47039 20404 47048
rect 20352 47005 20361 47039
rect 20361 47005 20395 47039
rect 20395 47005 20404 47039
rect 20352 46996 20404 47005
rect 32404 47064 32456 47116
rect 33232 47064 33284 47116
rect 43628 47107 43680 47116
rect 43628 47073 43637 47107
rect 43637 47073 43671 47107
rect 43671 47073 43680 47107
rect 43628 47064 43680 47073
rect 44732 47064 44784 47116
rect 46756 47107 46808 47116
rect 46756 47073 46765 47107
rect 46765 47073 46799 47107
rect 46799 47073 46808 47107
rect 46756 47064 46808 47073
rect 28264 46996 28316 47048
rect 42708 46996 42760 47048
rect 45008 47039 45060 47048
rect 45008 47005 45017 47039
rect 45017 47005 45051 47039
rect 45051 47005 45060 47039
rect 45008 46996 45060 47005
rect 45652 47039 45704 47048
rect 45652 47005 45661 47039
rect 45661 47005 45695 47039
rect 45695 47005 45704 47039
rect 45652 46996 45704 47005
rect 47952 46996 48004 47048
rect 48964 46996 49016 47048
rect 39304 46928 39356 46980
rect 41512 46928 41564 46980
rect 41788 46928 41840 46980
rect 42340 46971 42392 46980
rect 42340 46937 42349 46971
rect 42349 46937 42383 46971
rect 42383 46937 42392 46971
rect 42340 46928 42392 46937
rect 45836 46928 45888 46980
rect 45744 46903 45796 46912
rect 45744 46869 45753 46903
rect 45753 46869 45787 46903
rect 45787 46869 45796 46903
rect 45744 46860 45796 46869
rect 19574 46758 19626 46810
rect 19638 46758 19690 46810
rect 19702 46758 19754 46810
rect 19766 46758 19818 46810
rect 19830 46758 19882 46810
rect 2872 46699 2924 46708
rect 2872 46665 2881 46699
rect 2881 46665 2915 46699
rect 2915 46665 2924 46699
rect 2872 46656 2924 46665
rect 44088 46699 44140 46708
rect 44088 46665 44097 46699
rect 44097 46665 44131 46699
rect 44131 46665 44140 46699
rect 44088 46656 44140 46665
rect 1952 46520 2004 46572
rect 2044 46563 2096 46572
rect 2044 46529 2053 46563
rect 2053 46529 2087 46563
rect 2087 46529 2096 46563
rect 2044 46520 2096 46529
rect 2320 46520 2372 46572
rect 11520 46588 11572 46640
rect 23664 46588 23716 46640
rect 24768 46588 24820 46640
rect 3608 46563 3660 46572
rect 3608 46529 3617 46563
rect 3617 46529 3651 46563
rect 3651 46529 3660 46563
rect 3608 46520 3660 46529
rect 4712 46520 4764 46572
rect 5356 46563 5408 46572
rect 5356 46529 5365 46563
rect 5365 46529 5399 46563
rect 5399 46529 5408 46563
rect 5356 46520 5408 46529
rect 42708 46520 42760 46572
rect 45008 46588 45060 46640
rect 45744 46588 45796 46640
rect 47032 46631 47084 46640
rect 47032 46597 47041 46631
rect 47041 46597 47075 46631
rect 47075 46597 47084 46631
rect 47032 46588 47084 46597
rect 47952 46631 48004 46640
rect 47952 46597 47961 46631
rect 47961 46597 47995 46631
rect 47995 46597 48004 46631
rect 47952 46588 48004 46597
rect 42800 46495 42852 46504
rect 42800 46461 42809 46495
rect 42809 46461 42843 46495
rect 42843 46461 42852 46495
rect 42800 46452 42852 46461
rect 44180 46452 44232 46504
rect 1768 46316 1820 46368
rect 47768 46316 47820 46368
rect 4214 46214 4266 46266
rect 4278 46214 4330 46266
rect 4342 46214 4394 46266
rect 4406 46214 4458 46266
rect 4470 46214 4522 46266
rect 34934 46214 34986 46266
rect 34998 46214 35050 46266
rect 35062 46214 35114 46266
rect 35126 46214 35178 46266
rect 35190 46214 35242 46266
rect 1584 46112 1636 46164
rect 3884 46112 3936 46164
rect 42708 46112 42760 46164
rect 43996 46112 44048 46164
rect 44824 46112 44876 46164
rect 45376 46112 45428 46164
rect 46480 46112 46532 46164
rect 30564 46044 30616 46096
rect 31668 46044 31720 46096
rect 1400 45951 1452 45960
rect 1400 45917 1409 45951
rect 1409 45917 1443 45951
rect 1443 45917 1452 45951
rect 1400 45908 1452 45917
rect 2320 45951 2372 45960
rect 2320 45917 2329 45951
rect 2329 45917 2363 45951
rect 2363 45917 2372 45951
rect 2320 45908 2372 45917
rect 3148 45951 3200 45960
rect 3148 45917 3157 45951
rect 3157 45917 3191 45951
rect 3191 45917 3200 45951
rect 3148 45908 3200 45917
rect 21364 45772 21416 45824
rect 26424 45772 26476 45824
rect 44364 45908 44416 45960
rect 46756 45976 46808 46028
rect 48136 46019 48188 46028
rect 48136 45985 48145 46019
rect 48145 45985 48179 46019
rect 48179 45985 48188 46019
rect 48136 45976 48188 45985
rect 46296 45951 46348 45960
rect 46296 45917 46305 45951
rect 46305 45917 46339 45951
rect 46339 45917 46348 45951
rect 46296 45908 46348 45917
rect 47676 45840 47728 45892
rect 47216 45772 47268 45824
rect 19574 45670 19626 45722
rect 19638 45670 19690 45722
rect 19702 45670 19754 45722
rect 19766 45670 19818 45722
rect 19830 45670 19882 45722
rect 3148 45500 3200 45552
rect 28264 45500 28316 45552
rect 44180 45432 44232 45484
rect 44732 45475 44784 45484
rect 44732 45441 44741 45475
rect 44741 45441 44775 45475
rect 44775 45441 44784 45475
rect 44732 45432 44784 45441
rect 47676 45543 47728 45552
rect 47676 45509 47685 45543
rect 47685 45509 47719 45543
rect 47719 45509 47728 45543
rect 47676 45500 47728 45509
rect 1952 45407 2004 45416
rect 1952 45373 1961 45407
rect 1961 45373 1995 45407
rect 1995 45373 2004 45407
rect 1952 45364 2004 45373
rect 2780 45407 2832 45416
rect 2780 45373 2789 45407
rect 2789 45373 2823 45407
rect 2823 45373 2832 45407
rect 2780 45364 2832 45373
rect 45192 45407 45244 45416
rect 45192 45373 45201 45407
rect 45201 45373 45235 45407
rect 45235 45373 45244 45407
rect 45192 45364 45244 45373
rect 46848 45407 46900 45416
rect 46848 45373 46857 45407
rect 46857 45373 46891 45407
rect 46891 45373 46900 45407
rect 46848 45364 46900 45373
rect 47676 45296 47728 45348
rect 4214 45126 4266 45178
rect 4278 45126 4330 45178
rect 4342 45126 4394 45178
rect 4406 45126 4458 45178
rect 4470 45126 4522 45178
rect 34934 45126 34986 45178
rect 34998 45126 35050 45178
rect 35062 45126 35114 45178
rect 35126 45126 35178 45178
rect 35190 45126 35242 45178
rect 45192 45067 45244 45076
rect 45192 45033 45201 45067
rect 45201 45033 45235 45067
rect 45235 45033 45244 45067
rect 45192 45024 45244 45033
rect 45560 45024 45612 45076
rect 45836 45024 45888 45076
rect 2780 44931 2832 44940
rect 2780 44897 2789 44931
rect 2789 44897 2823 44931
rect 2823 44897 2832 44931
rect 2780 44888 2832 44897
rect 46756 44888 46808 44940
rect 48136 44931 48188 44940
rect 48136 44897 48145 44931
rect 48145 44897 48179 44931
rect 48179 44897 48188 44931
rect 48136 44888 48188 44897
rect 45928 44820 45980 44872
rect 3424 44752 3476 44804
rect 46940 44752 46992 44804
rect 2872 44684 2924 44736
rect 19574 44582 19626 44634
rect 19638 44582 19690 44634
rect 19702 44582 19754 44634
rect 19766 44582 19818 44634
rect 19830 44582 19882 44634
rect 1952 44480 2004 44532
rect 3424 44523 3476 44532
rect 3424 44489 3433 44523
rect 3433 44489 3467 44523
rect 3467 44489 3476 44523
rect 3424 44480 3476 44489
rect 46940 44523 46992 44532
rect 46940 44489 46949 44523
rect 46949 44489 46983 44523
rect 46983 44489 46992 44523
rect 46940 44480 46992 44489
rect 47676 44523 47728 44532
rect 47676 44489 47685 44523
rect 47685 44489 47719 44523
rect 47719 44489 47728 44523
rect 47676 44480 47728 44489
rect 1860 44387 1912 44396
rect 1860 44353 1869 44387
rect 1869 44353 1903 44387
rect 1903 44353 1912 44387
rect 1860 44344 1912 44353
rect 2228 44344 2280 44396
rect 3332 44387 3384 44396
rect 3332 44353 3341 44387
rect 3341 44353 3375 44387
rect 3375 44353 3384 44387
rect 3332 44344 3384 44353
rect 45100 44344 45152 44396
rect 46296 44344 46348 44396
rect 46572 44344 46624 44396
rect 47492 44344 47544 44396
rect 36544 44276 36596 44328
rect 45560 44276 45612 44328
rect 20352 44208 20404 44260
rect 20536 44208 20588 44260
rect 43444 44208 43496 44260
rect 46020 44208 46072 44260
rect 2136 44183 2188 44192
rect 2136 44149 2145 44183
rect 2145 44149 2179 44183
rect 2179 44149 2188 44183
rect 2136 44140 2188 44149
rect 45652 44140 45704 44192
rect 45928 44140 45980 44192
rect 4214 44038 4266 44090
rect 4278 44038 4330 44090
rect 4342 44038 4394 44090
rect 4406 44038 4458 44090
rect 4470 44038 4522 44090
rect 34934 44038 34986 44090
rect 34998 44038 35050 44090
rect 35062 44038 35114 44090
rect 35126 44038 35178 44090
rect 35190 44038 35242 44090
rect 2872 43979 2924 43988
rect 2872 43945 2881 43979
rect 2881 43945 2915 43979
rect 2915 43945 2924 43979
rect 2872 43936 2924 43945
rect 46756 43979 46808 43988
rect 46756 43945 46765 43979
rect 46765 43945 46799 43979
rect 46799 43945 46808 43979
rect 46756 43936 46808 43945
rect 46664 43868 46716 43920
rect 21916 43800 21968 43852
rect 7748 43732 7800 43784
rect 26700 43732 26752 43784
rect 1860 43707 1912 43716
rect 1860 43673 1869 43707
rect 1869 43673 1903 43707
rect 1903 43673 1912 43707
rect 1860 43664 1912 43673
rect 47860 43775 47912 43784
rect 47860 43741 47869 43775
rect 47869 43741 47903 43775
rect 47903 43741 47912 43775
rect 47860 43732 47912 43741
rect 47492 43664 47544 43716
rect 48228 43664 48280 43716
rect 1676 43596 1728 43648
rect 46940 43596 46992 43648
rect 19574 43494 19626 43546
rect 19638 43494 19690 43546
rect 19702 43494 19754 43546
rect 19766 43494 19818 43546
rect 19830 43494 19882 43546
rect 23388 43392 23440 43444
rect 47308 43392 47360 43444
rect 47952 43299 48004 43308
rect 47952 43265 47961 43299
rect 47961 43265 47995 43299
rect 47995 43265 48004 43299
rect 47952 43256 48004 43265
rect 47032 43095 47084 43104
rect 47032 43061 47041 43095
rect 47041 43061 47075 43095
rect 47075 43061 47084 43095
rect 47032 43052 47084 43061
rect 48044 43095 48096 43104
rect 48044 43061 48053 43095
rect 48053 43061 48087 43095
rect 48087 43061 48096 43095
rect 48044 43052 48096 43061
rect 4214 42950 4266 43002
rect 4278 42950 4330 43002
rect 4342 42950 4394 43002
rect 4406 42950 4458 43002
rect 4470 42950 4522 43002
rect 34934 42950 34986 43002
rect 34998 42950 35050 43002
rect 35062 42950 35114 43002
rect 35126 42950 35178 43002
rect 35190 42950 35242 43002
rect 47032 42712 47084 42764
rect 48136 42755 48188 42764
rect 48136 42721 48145 42755
rect 48145 42721 48179 42755
rect 48179 42721 48188 42755
rect 48136 42712 48188 42721
rect 46480 42619 46532 42628
rect 46480 42585 46489 42619
rect 46489 42585 46523 42619
rect 46523 42585 46532 42619
rect 46480 42576 46532 42585
rect 19574 42406 19626 42458
rect 19638 42406 19690 42458
rect 19702 42406 19754 42458
rect 19766 42406 19818 42458
rect 19830 42406 19882 42458
rect 45744 42236 45796 42288
rect 46480 42236 46532 42288
rect 22928 42211 22980 42220
rect 20720 42100 20772 42152
rect 22928 42177 22937 42211
rect 22937 42177 22971 42211
rect 22971 42177 22980 42211
rect 22928 42168 22980 42177
rect 24584 42168 24636 42220
rect 47216 42168 47268 42220
rect 47860 42211 47912 42220
rect 47860 42177 47869 42211
rect 47869 42177 47903 42211
rect 47903 42177 47912 42211
rect 47860 42168 47912 42177
rect 25872 42100 25924 42152
rect 1400 41964 1452 42016
rect 23572 41964 23624 42016
rect 4214 41862 4266 41914
rect 4278 41862 4330 41914
rect 4342 41862 4394 41914
rect 4406 41862 4458 41914
rect 4470 41862 4522 41914
rect 34934 41862 34986 41914
rect 34998 41862 35050 41914
rect 35062 41862 35114 41914
rect 35126 41862 35178 41914
rect 35190 41862 35242 41914
rect 1400 41667 1452 41676
rect 1400 41633 1409 41667
rect 1409 41633 1443 41667
rect 1443 41633 1452 41667
rect 1400 41624 1452 41633
rect 1860 41667 1912 41676
rect 1860 41633 1869 41667
rect 1869 41633 1903 41667
rect 1903 41633 1912 41667
rect 1860 41624 1912 41633
rect 19340 41556 19392 41608
rect 48044 41692 48096 41744
rect 47676 41624 47728 41676
rect 1584 41531 1636 41540
rect 1584 41497 1593 41531
rect 1593 41497 1627 41531
rect 1627 41497 1636 41531
rect 1584 41488 1636 41497
rect 19432 41420 19484 41472
rect 21824 41488 21876 41540
rect 22376 41488 22428 41540
rect 23020 41488 23072 41540
rect 23572 41599 23624 41608
rect 23572 41565 23581 41599
rect 23581 41565 23615 41599
rect 23615 41565 23624 41599
rect 23756 41599 23808 41608
rect 23572 41556 23624 41565
rect 23756 41565 23765 41599
rect 23765 41565 23799 41599
rect 23799 41565 23808 41599
rect 23756 41556 23808 41565
rect 46480 41531 46532 41540
rect 46480 41497 46489 41531
rect 46489 41497 46523 41531
rect 46523 41497 46532 41531
rect 46480 41488 46532 41497
rect 48136 41531 48188 41540
rect 48136 41497 48145 41531
rect 48145 41497 48179 41531
rect 48179 41497 48188 41531
rect 48136 41488 48188 41497
rect 20904 41420 20956 41472
rect 22192 41420 22244 41472
rect 23480 41420 23532 41472
rect 19574 41318 19626 41370
rect 19638 41318 19690 41370
rect 19702 41318 19754 41370
rect 19766 41318 19818 41370
rect 19830 41318 19882 41370
rect 1584 41216 1636 41268
rect 19432 41216 19484 41268
rect 21824 41259 21876 41268
rect 21824 41225 21833 41259
rect 21833 41225 21867 41259
rect 21867 41225 21876 41259
rect 21824 41216 21876 41225
rect 1860 41123 1912 41132
rect 1860 41089 1869 41123
rect 1869 41089 1903 41123
rect 1903 41089 1912 41123
rect 1860 41080 1912 41089
rect 2320 41080 2372 41132
rect 21916 41148 21968 41200
rect 2964 41080 3016 41132
rect 18788 41012 18840 41064
rect 20076 41080 20128 41132
rect 2412 40944 2464 40996
rect 20904 41080 20956 41132
rect 22284 41216 22336 41268
rect 46480 41216 46532 41268
rect 23480 41191 23532 41200
rect 23480 41157 23514 41191
rect 23514 41157 23532 41191
rect 23480 41148 23532 41157
rect 20812 41012 20864 41064
rect 22284 41123 22336 41132
rect 22284 41089 22293 41123
rect 22293 41089 22327 41123
rect 22327 41089 22336 41123
rect 22284 41080 22336 41089
rect 23756 41080 23808 41132
rect 46664 41123 46716 41132
rect 46664 41089 46673 41123
rect 46673 41089 46707 41123
rect 46707 41089 46716 41123
rect 46664 41080 46716 41089
rect 47676 41080 47728 41132
rect 22376 41012 22428 41064
rect 23204 41055 23256 41064
rect 23204 41021 23213 41055
rect 23213 41021 23247 41055
rect 23247 41021 23256 41055
rect 23204 41012 23256 41021
rect 19984 40876 20036 40928
rect 20720 40944 20772 40996
rect 24676 40876 24728 40928
rect 4214 40774 4266 40826
rect 4278 40774 4330 40826
rect 4342 40774 4394 40826
rect 4406 40774 4458 40826
rect 4470 40774 4522 40826
rect 34934 40774 34986 40826
rect 34998 40774 35050 40826
rect 35062 40774 35114 40826
rect 35126 40774 35178 40826
rect 35190 40774 35242 40826
rect 22284 40672 22336 40724
rect 1400 40511 1452 40520
rect 1400 40477 1409 40511
rect 1409 40477 1443 40511
rect 1443 40477 1452 40511
rect 1400 40468 1452 40477
rect 18604 40468 18656 40520
rect 20444 40468 20496 40520
rect 22100 40511 22152 40520
rect 22100 40477 22109 40511
rect 22109 40477 22143 40511
rect 22143 40477 22152 40511
rect 29828 40672 29880 40724
rect 22652 40536 22704 40588
rect 23204 40536 23256 40588
rect 47308 40579 47360 40588
rect 47308 40545 47317 40579
rect 47317 40545 47351 40579
rect 47351 40545 47360 40579
rect 47308 40536 47360 40545
rect 22100 40468 22152 40477
rect 22928 40511 22980 40520
rect 22928 40477 22937 40511
rect 22937 40477 22971 40511
rect 22971 40477 22980 40511
rect 22928 40468 22980 40477
rect 47400 40468 47452 40520
rect 23112 40400 23164 40452
rect 24584 40400 24636 40452
rect 24860 40400 24912 40452
rect 1584 40375 1636 40384
rect 1584 40341 1593 40375
rect 1593 40341 1627 40375
rect 1627 40341 1636 40375
rect 1584 40332 1636 40341
rect 19432 40375 19484 40384
rect 19432 40341 19441 40375
rect 19441 40341 19475 40375
rect 19475 40341 19484 40375
rect 19432 40332 19484 40341
rect 20812 40332 20864 40384
rect 22928 40332 22980 40384
rect 24492 40332 24544 40384
rect 19574 40230 19626 40282
rect 19638 40230 19690 40282
rect 19702 40230 19754 40282
rect 19766 40230 19818 40282
rect 19830 40230 19882 40282
rect 20444 40171 20496 40180
rect 20444 40137 20453 40171
rect 20453 40137 20487 40171
rect 20487 40137 20496 40171
rect 20444 40128 20496 40137
rect 22928 40128 22980 40180
rect 24584 40171 24636 40180
rect 24584 40137 24593 40171
rect 24593 40137 24627 40171
rect 24627 40137 24636 40171
rect 24584 40128 24636 40137
rect 26608 40128 26660 40180
rect 19892 40060 19944 40112
rect 20076 40060 20128 40112
rect 23756 40060 23808 40112
rect 18512 39992 18564 40044
rect 19156 39992 19208 40044
rect 22836 39992 22888 40044
rect 24124 39992 24176 40044
rect 25320 40060 25372 40112
rect 27344 40103 27396 40112
rect 25044 40035 25096 40044
rect 25044 40001 25053 40035
rect 25053 40001 25087 40035
rect 25087 40001 25096 40035
rect 25044 39992 25096 40001
rect 25872 40035 25924 40044
rect 18788 39856 18840 39908
rect 22192 39924 22244 39976
rect 22652 39924 22704 39976
rect 23848 39924 23900 39976
rect 25872 40001 25881 40035
rect 25881 40001 25915 40035
rect 25915 40001 25924 40035
rect 25872 39992 25924 40001
rect 27344 40069 27353 40103
rect 27353 40069 27387 40103
rect 27387 40069 27396 40103
rect 27344 40060 27396 40069
rect 25780 39924 25832 39976
rect 19340 39788 19392 39840
rect 20628 39856 20680 39908
rect 24952 39856 25004 39908
rect 27528 39967 27580 39976
rect 27528 39933 27537 39967
rect 27537 39933 27571 39967
rect 27571 39933 27580 39967
rect 28080 39992 28132 40044
rect 43628 39992 43680 40044
rect 47492 39992 47544 40044
rect 27528 39924 27580 39933
rect 29000 39924 29052 39976
rect 24860 39788 24912 39840
rect 26148 39788 26200 39840
rect 28908 39788 28960 39840
rect 46296 39788 46348 39840
rect 47676 39831 47728 39840
rect 47676 39797 47685 39831
rect 47685 39797 47719 39831
rect 47719 39797 47728 39831
rect 47676 39788 47728 39797
rect 4214 39686 4266 39738
rect 4278 39686 4330 39738
rect 4342 39686 4394 39738
rect 4406 39686 4458 39738
rect 4470 39686 4522 39738
rect 34934 39686 34986 39738
rect 34998 39686 35050 39738
rect 35062 39686 35114 39738
rect 35126 39686 35178 39738
rect 35190 39686 35242 39738
rect 19156 39584 19208 39636
rect 22836 39584 22888 39636
rect 19432 39448 19484 39500
rect 20812 39491 20864 39500
rect 19340 39380 19392 39432
rect 20812 39457 20821 39491
rect 20821 39457 20855 39491
rect 20855 39457 20864 39491
rect 20812 39448 20864 39457
rect 48044 39584 48096 39636
rect 28080 39516 28132 39568
rect 19892 39423 19944 39432
rect 17408 39312 17460 39364
rect 17224 39244 17276 39296
rect 18696 39287 18748 39296
rect 18696 39253 18705 39287
rect 18705 39253 18739 39287
rect 18739 39253 18748 39287
rect 18696 39244 18748 39253
rect 18788 39244 18840 39296
rect 19892 39389 19901 39423
rect 19901 39389 19935 39423
rect 19935 39389 19944 39423
rect 19892 39380 19944 39389
rect 20076 39380 20128 39432
rect 20720 39380 20772 39432
rect 26056 39448 26108 39500
rect 28448 39448 28500 39500
rect 23112 39423 23164 39432
rect 23112 39389 23121 39423
rect 23121 39389 23155 39423
rect 23155 39389 23164 39423
rect 23112 39380 23164 39389
rect 23848 39380 23900 39432
rect 24492 39380 24544 39432
rect 28540 39380 28592 39432
rect 23756 39312 23808 39364
rect 23020 39244 23072 39296
rect 24032 39244 24084 39296
rect 24676 39312 24728 39364
rect 25688 39312 25740 39364
rect 25136 39244 25188 39296
rect 25780 39244 25832 39296
rect 27804 39244 27856 39296
rect 28356 39287 28408 39296
rect 28356 39253 28365 39287
rect 28365 39253 28399 39287
rect 28399 39253 28408 39287
rect 28356 39244 28408 39253
rect 29000 39423 29052 39432
rect 29000 39389 29009 39423
rect 29009 39389 29043 39423
rect 29043 39389 29052 39423
rect 46296 39491 46348 39500
rect 46296 39457 46305 39491
rect 46305 39457 46339 39491
rect 46339 39457 46348 39491
rect 46296 39448 46348 39457
rect 47676 39448 47728 39500
rect 48136 39491 48188 39500
rect 48136 39457 48145 39491
rect 48145 39457 48179 39491
rect 48179 39457 48188 39491
rect 48136 39448 48188 39457
rect 29000 39380 29052 39389
rect 28908 39312 28960 39364
rect 28816 39244 28868 39296
rect 29828 39244 29880 39296
rect 19574 39142 19626 39194
rect 19638 39142 19690 39194
rect 19702 39142 19754 39194
rect 19766 39142 19818 39194
rect 19830 39142 19882 39194
rect 17408 39083 17460 39092
rect 17408 39049 17417 39083
rect 17417 39049 17451 39083
rect 17451 39049 17460 39083
rect 17408 39040 17460 39049
rect 20720 39040 20772 39092
rect 23848 39040 23900 39092
rect 25044 39040 25096 39092
rect 25688 39083 25740 39092
rect 25688 39049 25697 39083
rect 25697 39049 25731 39083
rect 25731 39049 25740 39083
rect 25688 39040 25740 39049
rect 27804 39083 27856 39092
rect 27804 39049 27813 39083
rect 27813 39049 27847 39083
rect 27847 39049 27856 39083
rect 27804 39040 27856 39049
rect 17592 38904 17644 38956
rect 19708 38972 19760 39024
rect 24032 39015 24084 39024
rect 24032 38981 24041 39015
rect 24041 38981 24075 39015
rect 24075 38981 24084 39015
rect 24032 38972 24084 38981
rect 18512 38947 18564 38956
rect 2044 38879 2096 38888
rect 2044 38845 2053 38879
rect 2053 38845 2087 38879
rect 2087 38845 2096 38879
rect 2044 38836 2096 38845
rect 2780 38836 2832 38888
rect 2872 38879 2924 38888
rect 2872 38845 2881 38879
rect 2881 38845 2915 38879
rect 2915 38845 2924 38879
rect 2872 38836 2924 38845
rect 17868 38768 17920 38820
rect 18512 38913 18521 38947
rect 18521 38913 18555 38947
rect 18555 38913 18564 38947
rect 18512 38904 18564 38913
rect 19800 38904 19852 38956
rect 24952 38972 25004 39024
rect 25136 38972 25188 39024
rect 18696 38836 18748 38888
rect 24216 38947 24268 38956
rect 24216 38913 24225 38947
rect 24225 38913 24259 38947
rect 24259 38913 24268 38947
rect 24216 38904 24268 38913
rect 25780 38904 25832 38956
rect 22284 38836 22336 38888
rect 25228 38836 25280 38888
rect 26148 38947 26200 38956
rect 26148 38913 26157 38947
rect 26157 38913 26191 38947
rect 26191 38913 26200 38947
rect 27344 38972 27396 39024
rect 48044 39083 48096 39092
rect 48044 39049 48053 39083
rect 48053 39049 48087 39083
rect 48087 39049 48096 39083
rect 48044 39040 48096 39049
rect 28356 38972 28408 39024
rect 26148 38904 26200 38913
rect 27804 38904 27856 38956
rect 28540 38947 28592 38956
rect 28540 38913 28549 38947
rect 28549 38913 28583 38947
rect 28583 38913 28592 38947
rect 28540 38904 28592 38913
rect 47952 38947 48004 38956
rect 47952 38913 47961 38947
rect 47961 38913 47995 38947
rect 47995 38913 48004 38947
rect 47952 38904 48004 38913
rect 18788 38700 18840 38752
rect 24952 38743 25004 38752
rect 24952 38709 24961 38743
rect 24961 38709 24995 38743
rect 24995 38709 25004 38743
rect 24952 38700 25004 38709
rect 25136 38700 25188 38752
rect 26056 38700 26108 38752
rect 27528 38836 27580 38888
rect 27344 38743 27396 38752
rect 27344 38709 27353 38743
rect 27353 38709 27387 38743
rect 27387 38709 27396 38743
rect 27344 38700 27396 38709
rect 47032 38743 47084 38752
rect 47032 38709 47041 38743
rect 47041 38709 47075 38743
rect 47075 38709 47084 38743
rect 47032 38700 47084 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 2044 38496 2096 38548
rect 21272 38496 21324 38548
rect 22928 38496 22980 38548
rect 27804 38496 27856 38548
rect 17868 38428 17920 38480
rect 20076 38428 20128 38480
rect 18420 38360 18472 38412
rect 25320 38428 25372 38480
rect 28540 38428 28592 38480
rect 22100 38360 22152 38412
rect 23112 38360 23164 38412
rect 24216 38360 24268 38412
rect 21088 38292 21140 38344
rect 22376 38335 22428 38344
rect 22376 38301 22385 38335
rect 22385 38301 22419 38335
rect 22419 38301 22428 38335
rect 22376 38292 22428 38301
rect 17040 38224 17092 38276
rect 18512 38224 18564 38276
rect 19340 38224 19392 38276
rect 19708 38267 19760 38276
rect 19708 38233 19717 38267
rect 19717 38233 19751 38267
rect 19751 38233 19760 38267
rect 19708 38224 19760 38233
rect 22836 38292 22888 38344
rect 23572 38292 23624 38344
rect 24952 38335 25004 38344
rect 24952 38301 24961 38335
rect 24961 38301 24995 38335
rect 24995 38301 25004 38335
rect 24952 38292 25004 38301
rect 25136 38335 25188 38344
rect 25136 38301 25145 38335
rect 25145 38301 25179 38335
rect 25179 38301 25188 38335
rect 25136 38292 25188 38301
rect 27344 38292 27396 38344
rect 28080 38360 28132 38412
rect 28448 38360 28500 38412
rect 28632 38335 28684 38344
rect 28632 38301 28641 38335
rect 28641 38301 28675 38335
rect 28675 38301 28684 38335
rect 28632 38292 28684 38301
rect 47032 38360 47084 38412
rect 48228 38360 48280 38412
rect 28908 38292 28960 38344
rect 29092 38292 29144 38344
rect 23020 38224 23072 38276
rect 24676 38224 24728 38276
rect 46940 38224 46992 38276
rect 18420 38199 18472 38208
rect 18420 38165 18429 38199
rect 18429 38165 18463 38199
rect 18463 38165 18472 38199
rect 18420 38156 18472 38165
rect 22008 38199 22060 38208
rect 22008 38165 22017 38199
rect 22017 38165 22051 38199
rect 22051 38165 22060 38199
rect 22008 38156 22060 38165
rect 25688 38156 25740 38208
rect 28908 38156 28960 38208
rect 19574 38054 19626 38106
rect 19638 38054 19690 38106
rect 19702 38054 19754 38106
rect 19766 38054 19818 38106
rect 19830 38054 19882 38106
rect 2780 37952 2832 38004
rect 24860 37952 24912 38004
rect 24952 37952 25004 38004
rect 46940 37995 46992 38004
rect 46940 37961 46949 37995
rect 46949 37961 46983 37995
rect 46983 37961 46992 37995
rect 46940 37952 46992 37961
rect 17132 37884 17184 37936
rect 1860 37859 1912 37868
rect 1860 37825 1869 37859
rect 1869 37825 1903 37859
rect 1903 37825 1912 37859
rect 1860 37816 1912 37825
rect 7288 37816 7340 37868
rect 18328 37816 18380 37868
rect 19432 37816 19484 37868
rect 22008 37884 22060 37936
rect 22836 37884 22888 37936
rect 22376 37816 22428 37868
rect 25136 37816 25188 37868
rect 21180 37748 21232 37800
rect 22192 37748 22244 37800
rect 24952 37791 25004 37800
rect 24952 37757 24961 37791
rect 24961 37757 24995 37791
rect 24995 37757 25004 37791
rect 24952 37748 25004 37757
rect 29000 37884 29052 37936
rect 25780 37859 25832 37868
rect 25780 37825 25789 37859
rect 25789 37825 25823 37859
rect 25823 37825 25832 37859
rect 25780 37816 25832 37825
rect 29184 37859 29236 37868
rect 29184 37825 29193 37859
rect 29193 37825 29227 37859
rect 29227 37825 29236 37859
rect 29184 37816 29236 37825
rect 27804 37748 27856 37800
rect 20996 37680 21048 37732
rect 25320 37680 25372 37732
rect 28448 37680 28500 37732
rect 29368 37859 29420 37868
rect 29368 37825 29377 37859
rect 29377 37825 29411 37859
rect 29411 37825 29420 37859
rect 29368 37816 29420 37825
rect 47308 37816 47360 37868
rect 47860 37859 47912 37868
rect 47860 37825 47869 37859
rect 47869 37825 47903 37859
rect 47903 37825 47912 37859
rect 47860 37816 47912 37825
rect 1952 37655 2004 37664
rect 1952 37621 1961 37655
rect 1961 37621 1995 37655
rect 1995 37621 2004 37655
rect 1952 37612 2004 37621
rect 18604 37655 18656 37664
rect 18604 37621 18613 37655
rect 18613 37621 18647 37655
rect 18647 37621 18656 37655
rect 18604 37612 18656 37621
rect 21088 37612 21140 37664
rect 24308 37655 24360 37664
rect 24308 37621 24317 37655
rect 24317 37621 24351 37655
rect 24351 37621 24360 37655
rect 24308 37612 24360 37621
rect 26240 37612 26292 37664
rect 27252 37612 27304 37664
rect 29644 37612 29696 37664
rect 48044 37655 48096 37664
rect 48044 37621 48053 37655
rect 48053 37621 48087 37655
rect 48087 37621 48096 37655
rect 48044 37612 48096 37621
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 1952 37408 2004 37460
rect 18328 37408 18380 37460
rect 23020 37408 23072 37460
rect 19156 37340 19208 37392
rect 1400 37315 1452 37324
rect 1400 37281 1409 37315
rect 1409 37281 1443 37315
rect 1443 37281 1452 37315
rect 1400 37272 1452 37281
rect 4068 37272 4120 37324
rect 8300 37272 8352 37324
rect 19064 37272 19116 37324
rect 19340 37272 19392 37324
rect 19984 37272 20036 37324
rect 22744 37272 22796 37324
rect 26240 37340 26292 37392
rect 27804 37340 27856 37392
rect 28540 37340 28592 37392
rect 7288 37247 7340 37256
rect 2136 37136 2188 37188
rect 2320 37136 2372 37188
rect 7288 37213 7297 37247
rect 7297 37213 7331 37247
rect 7331 37213 7340 37247
rect 7288 37204 7340 37213
rect 16488 37204 16540 37256
rect 20444 37204 20496 37256
rect 20628 37204 20680 37256
rect 21088 37204 21140 37256
rect 24308 37204 24360 37256
rect 24952 37272 25004 37324
rect 26148 37272 26200 37324
rect 33048 37272 33100 37324
rect 46848 37272 46900 37324
rect 29644 37204 29696 37256
rect 46296 37247 46348 37256
rect 46296 37213 46305 37247
rect 46305 37213 46339 37247
rect 46339 37213 46348 37247
rect 46296 37204 46348 37213
rect 17224 37136 17276 37188
rect 17684 37136 17736 37188
rect 7380 37111 7432 37120
rect 7380 37077 7389 37111
rect 7389 37077 7423 37111
rect 7423 37077 7432 37111
rect 7380 37068 7432 37077
rect 22744 37068 22796 37120
rect 23756 37136 23808 37188
rect 25780 37136 25832 37188
rect 27068 37136 27120 37188
rect 47676 37136 47728 37188
rect 48136 37179 48188 37188
rect 48136 37145 48145 37179
rect 48145 37145 48179 37179
rect 48179 37145 48188 37179
rect 48136 37136 48188 37145
rect 24400 37111 24452 37120
rect 24400 37077 24409 37111
rect 24409 37077 24443 37111
rect 24443 37077 24452 37111
rect 24400 37068 24452 37077
rect 25872 37068 25924 37120
rect 29644 37068 29696 37120
rect 30932 37111 30984 37120
rect 30932 37077 30941 37111
rect 30941 37077 30975 37111
rect 30975 37077 30984 37111
rect 30932 37068 30984 37077
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 21180 36864 21232 36916
rect 25780 36907 25832 36916
rect 25780 36873 25789 36907
rect 25789 36873 25823 36907
rect 25823 36873 25832 36907
rect 25780 36864 25832 36873
rect 29368 36864 29420 36916
rect 47676 36907 47728 36916
rect 47676 36873 47685 36907
rect 47685 36873 47719 36907
rect 47719 36873 47728 36907
rect 47676 36864 47728 36873
rect 7380 36839 7432 36848
rect 7380 36805 7389 36839
rect 7389 36805 7423 36839
rect 7423 36805 7432 36839
rect 7380 36796 7432 36805
rect 17408 36796 17460 36848
rect 24400 36796 24452 36848
rect 24584 36796 24636 36848
rect 46388 36796 46440 36848
rect 18052 36771 18104 36780
rect 18052 36737 18061 36771
rect 18061 36737 18095 36771
rect 18095 36737 18104 36771
rect 18052 36728 18104 36737
rect 8208 36660 8260 36712
rect 8300 36703 8352 36712
rect 8300 36669 8309 36703
rect 8309 36669 8343 36703
rect 8343 36669 8352 36703
rect 8300 36660 8352 36669
rect 17132 36592 17184 36644
rect 18052 36592 18104 36644
rect 18236 36771 18288 36780
rect 18236 36737 18245 36771
rect 18245 36737 18279 36771
rect 18279 36737 18288 36771
rect 18236 36728 18288 36737
rect 18328 36660 18380 36712
rect 19340 36728 19392 36780
rect 23572 36728 23624 36780
rect 23756 36728 23808 36780
rect 25872 36728 25924 36780
rect 26976 36728 27028 36780
rect 27804 36771 27856 36780
rect 27804 36737 27813 36771
rect 27813 36737 27847 36771
rect 27847 36737 27856 36771
rect 27804 36728 27856 36737
rect 27896 36728 27948 36780
rect 29828 36771 29880 36780
rect 29828 36737 29837 36771
rect 29837 36737 29871 36771
rect 29871 36737 29880 36771
rect 29828 36728 29880 36737
rect 30012 36771 30064 36780
rect 30012 36737 30021 36771
rect 30021 36737 30055 36771
rect 30055 36737 30064 36771
rect 30012 36728 30064 36737
rect 19892 36703 19944 36712
rect 19892 36669 19901 36703
rect 19901 36669 19935 36703
rect 19935 36669 19944 36703
rect 19892 36660 19944 36669
rect 20996 36660 21048 36712
rect 26148 36660 26200 36712
rect 30932 36728 30984 36780
rect 46296 36728 46348 36780
rect 20628 36592 20680 36644
rect 23572 36592 23624 36644
rect 2044 36524 2096 36576
rect 18144 36524 18196 36576
rect 19248 36567 19300 36576
rect 19248 36533 19257 36567
rect 19257 36533 19291 36567
rect 19291 36533 19300 36567
rect 19248 36524 19300 36533
rect 20904 36524 20956 36576
rect 24584 36524 24636 36576
rect 25964 36524 26016 36576
rect 26332 36524 26384 36576
rect 27068 36524 27120 36576
rect 29644 36524 29696 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 3332 36320 3384 36372
rect 8208 36363 8260 36372
rect 8208 36329 8217 36363
rect 8217 36329 8251 36363
rect 8251 36329 8260 36363
rect 8208 36320 8260 36329
rect 17132 36363 17184 36372
rect 17132 36329 17141 36363
rect 17141 36329 17175 36363
rect 17175 36329 17184 36363
rect 17132 36320 17184 36329
rect 17684 36363 17736 36372
rect 17684 36329 17693 36363
rect 17693 36329 17727 36363
rect 17727 36329 17736 36363
rect 17684 36320 17736 36329
rect 18236 36320 18288 36372
rect 19892 36320 19944 36372
rect 3332 36116 3384 36168
rect 15568 36116 15620 36168
rect 17040 36159 17092 36168
rect 17040 36125 17049 36159
rect 17049 36125 17083 36159
rect 17083 36125 17092 36159
rect 17040 36116 17092 36125
rect 17684 36116 17736 36168
rect 18604 36184 18656 36236
rect 20076 36252 20128 36304
rect 20444 36252 20496 36304
rect 18328 36159 18380 36168
rect 18328 36125 18337 36159
rect 18337 36125 18371 36159
rect 18371 36125 18380 36159
rect 18328 36116 18380 36125
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 19432 36159 19484 36168
rect 19432 36125 19441 36159
rect 19441 36125 19475 36159
rect 19475 36125 19484 36159
rect 19432 36116 19484 36125
rect 20904 36184 20956 36236
rect 22192 36320 22244 36372
rect 27896 36320 27948 36372
rect 22468 36252 22520 36304
rect 26792 36252 26844 36304
rect 23112 36116 23164 36168
rect 7656 36048 7708 36100
rect 3056 36023 3108 36032
rect 3056 35989 3065 36023
rect 3065 35989 3099 36023
rect 3099 35989 3108 36023
rect 3056 35980 3108 35989
rect 26332 36116 26384 36168
rect 28172 36252 28224 36304
rect 30012 36252 30064 36304
rect 27528 36159 27580 36168
rect 24400 36048 24452 36100
rect 25964 36091 26016 36100
rect 25964 36057 25973 36091
rect 25973 36057 26007 36091
rect 26007 36057 26016 36091
rect 25964 36048 26016 36057
rect 18512 35980 18564 36032
rect 20076 35980 20128 36032
rect 21088 35980 21140 36032
rect 23112 35980 23164 36032
rect 23204 35980 23256 36032
rect 24584 35980 24636 36032
rect 26884 36048 26936 36100
rect 27528 36125 27537 36159
rect 27537 36125 27571 36159
rect 27571 36125 27580 36159
rect 27528 36116 27580 36125
rect 47860 36159 47912 36168
rect 47860 36125 47869 36159
rect 47869 36125 47903 36159
rect 47903 36125 47912 36159
rect 47860 36116 47912 36125
rect 48136 35980 48188 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 1584 35776 1636 35828
rect 7656 35819 7708 35828
rect 3056 35708 3108 35760
rect 7656 35785 7665 35819
rect 7665 35785 7699 35819
rect 7699 35785 7708 35819
rect 7656 35776 7708 35785
rect 8392 35776 8444 35828
rect 24676 35776 24728 35828
rect 17408 35751 17460 35760
rect 2044 35683 2096 35692
rect 2044 35649 2053 35683
rect 2053 35649 2087 35683
rect 2087 35649 2096 35683
rect 2044 35640 2096 35649
rect 2780 35615 2832 35624
rect 2780 35581 2789 35615
rect 2789 35581 2823 35615
rect 2823 35581 2832 35615
rect 2780 35572 2832 35581
rect 17408 35717 17417 35751
rect 17417 35717 17451 35751
rect 17451 35717 17460 35751
rect 17408 35708 17460 35717
rect 18328 35708 18380 35760
rect 19892 35708 19944 35760
rect 20720 35708 20772 35760
rect 17960 35640 18012 35692
rect 18144 35683 18196 35692
rect 18144 35649 18178 35683
rect 18178 35649 18196 35683
rect 18144 35640 18196 35649
rect 20812 35640 20864 35692
rect 20996 35683 21048 35692
rect 20996 35649 21020 35683
rect 21020 35649 21048 35683
rect 20996 35640 21048 35649
rect 21088 35683 21140 35692
rect 21088 35649 21097 35683
rect 21097 35649 21131 35683
rect 21131 35649 21140 35683
rect 21088 35640 21140 35649
rect 21456 35640 21508 35692
rect 22192 35708 22244 35760
rect 24216 35708 24268 35760
rect 25780 35776 25832 35828
rect 21916 35640 21968 35692
rect 23664 35640 23716 35692
rect 24492 35640 24544 35692
rect 27804 35708 27856 35760
rect 15568 35572 15620 35624
rect 16488 35572 16540 35624
rect 23756 35572 23808 35624
rect 24584 35572 24636 35624
rect 27436 35640 27488 35692
rect 48228 35640 48280 35692
rect 26240 35615 26292 35624
rect 26240 35581 26249 35615
rect 26249 35581 26283 35615
rect 26283 35581 26292 35615
rect 26240 35572 26292 35581
rect 17132 35436 17184 35488
rect 19340 35436 19392 35488
rect 19800 35436 19852 35488
rect 27344 35504 27396 35556
rect 23296 35436 23348 35488
rect 27252 35436 27304 35488
rect 47216 35436 47268 35488
rect 48228 35436 48280 35488
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 15568 35275 15620 35284
rect 15568 35241 15577 35275
rect 15577 35241 15611 35275
rect 15611 35241 15620 35275
rect 15568 35232 15620 35241
rect 24584 35275 24636 35284
rect 13084 35096 13136 35148
rect 13268 35139 13320 35148
rect 13268 35105 13277 35139
rect 13277 35105 13311 35139
rect 13311 35105 13320 35139
rect 13268 35096 13320 35105
rect 1400 35071 1452 35080
rect 1400 35037 1409 35071
rect 1409 35037 1443 35071
rect 1443 35037 1452 35071
rect 1400 35028 1452 35037
rect 17408 35028 17460 35080
rect 17684 35164 17736 35216
rect 18972 35164 19024 35216
rect 19984 35096 20036 35148
rect 24584 35241 24593 35275
rect 24593 35241 24627 35275
rect 24627 35241 24636 35275
rect 24584 35232 24636 35241
rect 27436 35232 27488 35284
rect 27620 35232 27672 35284
rect 18049 35071 18101 35080
rect 18049 35037 18058 35071
rect 18058 35037 18092 35071
rect 18092 35037 18101 35071
rect 18049 35028 18101 35037
rect 18144 35071 18196 35080
rect 18144 35037 18158 35071
rect 18158 35037 18192 35071
rect 18192 35037 18196 35071
rect 18328 35071 18380 35080
rect 18144 35028 18196 35037
rect 18328 35037 18337 35071
rect 18337 35037 18371 35071
rect 18371 35037 18380 35071
rect 18328 35028 18380 35037
rect 19340 35028 19392 35080
rect 19616 35071 19668 35080
rect 19616 35037 19625 35071
rect 19625 35037 19659 35071
rect 19659 35037 19668 35071
rect 19616 35028 19668 35037
rect 21272 35096 21324 35148
rect 21548 35071 21600 35080
rect 11612 35003 11664 35012
rect 11612 34969 11621 35003
rect 11621 34969 11655 35003
rect 11655 34969 11664 35003
rect 11612 34960 11664 34969
rect 21548 35037 21571 35071
rect 21571 35037 21600 35071
rect 21548 35028 21600 35037
rect 24676 35164 24728 35216
rect 23204 35139 23256 35148
rect 23204 35105 23213 35139
rect 23213 35105 23247 35139
rect 23247 35105 23256 35139
rect 23204 35096 23256 35105
rect 23296 35096 23348 35148
rect 25504 35139 25556 35148
rect 25504 35105 25513 35139
rect 25513 35105 25547 35139
rect 25547 35105 25556 35139
rect 25504 35096 25556 35105
rect 25688 35139 25740 35148
rect 25688 35105 25697 35139
rect 25697 35105 25731 35139
rect 25731 35105 25740 35139
rect 25688 35096 25740 35105
rect 26792 35096 26844 35148
rect 21916 35071 21968 35080
rect 20720 34960 20772 35012
rect 20996 34960 21048 35012
rect 21916 35037 21925 35071
rect 21925 35037 21959 35071
rect 21959 35037 21968 35071
rect 21916 35028 21968 35037
rect 22008 35028 22060 35080
rect 26240 35028 26292 35080
rect 47032 35096 47084 35148
rect 48136 35139 48188 35148
rect 48136 35105 48145 35139
rect 48145 35105 48179 35139
rect 48179 35105 48188 35139
rect 48136 35096 48188 35105
rect 23480 34960 23532 35012
rect 24492 34960 24544 35012
rect 17684 34935 17736 34944
rect 17684 34901 17693 34935
rect 17693 34901 17727 34935
rect 17727 34901 17736 34935
rect 17684 34892 17736 34901
rect 19248 34935 19300 34944
rect 19248 34901 19257 34935
rect 19257 34901 19291 34935
rect 19291 34901 19300 34935
rect 19248 34892 19300 34901
rect 21916 34892 21968 34944
rect 25136 34960 25188 35012
rect 25596 34892 25648 34944
rect 27252 35071 27304 35080
rect 27252 35037 27261 35071
rect 27261 35037 27295 35071
rect 27295 35037 27304 35071
rect 27252 35028 27304 35037
rect 27528 35028 27580 35080
rect 32312 35071 32364 35080
rect 32312 35037 32321 35071
rect 32321 35037 32355 35071
rect 32355 35037 32364 35071
rect 32312 35028 32364 35037
rect 27988 35003 28040 35012
rect 27988 34969 27997 35003
rect 27997 34969 28031 35003
rect 28031 34969 28040 35003
rect 27988 34960 28040 34969
rect 33416 34960 33468 35012
rect 46480 35003 46532 35012
rect 46480 34969 46489 35003
rect 46489 34969 46523 35003
rect 46523 34969 46532 35003
rect 46480 34960 46532 34969
rect 27528 34892 27580 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 11612 34731 11664 34740
rect 11612 34697 11621 34731
rect 11621 34697 11655 34731
rect 11655 34697 11664 34731
rect 11612 34688 11664 34697
rect 19340 34688 19392 34740
rect 19432 34688 19484 34740
rect 20720 34688 20772 34740
rect 17684 34620 17736 34672
rect 22836 34688 22888 34740
rect 11520 34595 11572 34604
rect 11520 34561 11529 34595
rect 11529 34561 11563 34595
rect 11563 34561 11572 34595
rect 11520 34552 11572 34561
rect 11980 34552 12032 34604
rect 15568 34552 15620 34604
rect 19340 34552 19392 34604
rect 22192 34620 22244 34672
rect 24584 34688 24636 34740
rect 26608 34688 26660 34740
rect 32312 34688 32364 34740
rect 23480 34620 23532 34672
rect 24676 34620 24728 34672
rect 21272 34527 21324 34536
rect 21272 34493 21281 34527
rect 21281 34493 21315 34527
rect 21315 34493 21324 34527
rect 21272 34484 21324 34493
rect 21916 34552 21968 34604
rect 25320 34595 25372 34604
rect 25320 34561 25329 34595
rect 25329 34561 25363 34595
rect 25363 34561 25372 34595
rect 25320 34552 25372 34561
rect 26608 34552 26660 34604
rect 27344 34620 27396 34672
rect 28080 34552 28132 34604
rect 29000 34620 29052 34672
rect 29460 34595 29512 34604
rect 29460 34561 29469 34595
rect 29469 34561 29503 34595
rect 29503 34561 29512 34595
rect 29460 34552 29512 34561
rect 43444 34620 43496 34672
rect 29736 34595 29788 34604
rect 29736 34561 29745 34595
rect 29745 34561 29779 34595
rect 29779 34561 29788 34595
rect 29736 34552 29788 34561
rect 30104 34552 30156 34604
rect 31760 34552 31812 34604
rect 47308 34552 47360 34604
rect 23664 34527 23716 34536
rect 15200 34416 15252 34468
rect 16396 34416 16448 34468
rect 1400 34348 1452 34400
rect 23664 34493 23673 34527
rect 23673 34493 23707 34527
rect 23707 34493 23716 34527
rect 23664 34484 23716 34493
rect 23756 34484 23808 34536
rect 26148 34484 26200 34536
rect 30380 34484 30432 34536
rect 31944 34484 31996 34536
rect 32128 34527 32180 34536
rect 32128 34493 32137 34527
rect 32137 34493 32171 34527
rect 32171 34493 32180 34527
rect 32128 34484 32180 34493
rect 33876 34484 33928 34536
rect 34520 34527 34572 34536
rect 34520 34493 34529 34527
rect 34529 34493 34563 34527
rect 34563 34493 34572 34527
rect 34520 34484 34572 34493
rect 27804 34416 27856 34468
rect 28172 34416 28224 34468
rect 47032 34459 47084 34468
rect 47032 34425 47041 34459
rect 47041 34425 47075 34459
rect 47075 34425 47084 34459
rect 47032 34416 47084 34425
rect 23480 34348 23532 34400
rect 25136 34348 25188 34400
rect 25872 34348 25924 34400
rect 28080 34348 28132 34400
rect 28356 34348 28408 34400
rect 29184 34348 29236 34400
rect 33508 34348 33560 34400
rect 46296 34348 46348 34400
rect 47676 34391 47728 34400
rect 47676 34357 47685 34391
rect 47685 34357 47719 34391
rect 47719 34357 47728 34391
rect 47676 34348 47728 34357
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 13084 34144 13136 34196
rect 1400 34051 1452 34060
rect 1400 34017 1409 34051
rect 1409 34017 1443 34051
rect 1443 34017 1452 34051
rect 1400 34008 1452 34017
rect 2780 34051 2832 34060
rect 2780 34017 2789 34051
rect 2789 34017 2823 34051
rect 2823 34017 2832 34051
rect 2780 34008 2832 34017
rect 15568 33940 15620 33992
rect 18144 34144 18196 34196
rect 22744 34144 22796 34196
rect 25504 34144 25556 34196
rect 25964 34187 26016 34196
rect 25964 34153 25973 34187
rect 25973 34153 26007 34187
rect 26007 34153 26016 34187
rect 25964 34144 26016 34153
rect 26240 34187 26292 34196
rect 26240 34153 26249 34187
rect 26249 34153 26283 34187
rect 26283 34153 26292 34187
rect 26240 34144 26292 34153
rect 28080 34144 28132 34196
rect 31208 34144 31260 34196
rect 31760 34144 31812 34196
rect 34520 34144 34572 34196
rect 16396 34076 16448 34128
rect 23940 34076 23992 34128
rect 26976 34119 27028 34128
rect 26976 34085 26985 34119
rect 26985 34085 27019 34119
rect 27019 34085 27028 34119
rect 26976 34076 27028 34085
rect 21272 34008 21324 34060
rect 24860 34051 24912 34060
rect 19248 33940 19300 33992
rect 2136 33872 2188 33924
rect 15476 33872 15528 33924
rect 17500 33872 17552 33924
rect 19432 33872 19484 33924
rect 21824 33940 21876 33992
rect 24860 34017 24869 34051
rect 24869 34017 24903 34051
rect 24903 34017 24912 34051
rect 24860 34008 24912 34017
rect 22284 33872 22336 33924
rect 23480 33915 23532 33924
rect 23480 33881 23489 33915
rect 23489 33881 23523 33915
rect 23523 33881 23532 33915
rect 23480 33872 23532 33881
rect 23756 33872 23808 33924
rect 24676 33872 24728 33924
rect 25136 33940 25188 33992
rect 26332 34008 26384 34060
rect 26608 34008 26660 34060
rect 17040 33847 17092 33856
rect 17040 33813 17049 33847
rect 17049 33813 17083 33847
rect 17083 33813 17092 33847
rect 17040 33804 17092 33813
rect 17132 33804 17184 33856
rect 23572 33804 23624 33856
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 24400 33804 24452 33856
rect 27988 33940 28040 33992
rect 28356 33940 28408 33992
rect 29552 33983 29604 33992
rect 29552 33949 29561 33983
rect 29561 33949 29595 33983
rect 29595 33949 29604 33983
rect 29552 33940 29604 33949
rect 28632 33915 28684 33924
rect 28632 33881 28641 33915
rect 28641 33881 28675 33915
rect 28675 33881 28684 33915
rect 28632 33872 28684 33881
rect 29092 33872 29144 33924
rect 31208 33940 31260 33992
rect 32404 34008 32456 34060
rect 47216 34076 47268 34128
rect 47676 34008 47728 34060
rect 48136 34051 48188 34060
rect 48136 34017 48145 34051
rect 48145 34017 48179 34051
rect 48179 34017 48188 34051
rect 48136 34008 48188 34017
rect 31944 33940 31996 33992
rect 32128 33872 32180 33924
rect 33324 33940 33376 33992
rect 33968 33940 34020 33992
rect 32588 33872 32640 33924
rect 29000 33847 29052 33856
rect 29000 33813 29009 33847
rect 29009 33813 29043 33847
rect 29043 33813 29052 33847
rect 29000 33804 29052 33813
rect 30932 33847 30984 33856
rect 30932 33813 30941 33847
rect 30941 33813 30975 33847
rect 30975 33813 30984 33847
rect 30932 33804 30984 33813
rect 31760 33804 31812 33856
rect 33876 33847 33928 33856
rect 33876 33813 33885 33847
rect 33885 33813 33919 33847
rect 33919 33813 33928 33847
rect 33876 33804 33928 33813
rect 47952 33804 48004 33856
rect 48136 33804 48188 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 2136 33643 2188 33652
rect 2136 33609 2145 33643
rect 2145 33609 2179 33643
rect 2179 33609 2188 33643
rect 2136 33600 2188 33609
rect 15476 33643 15528 33652
rect 15476 33609 15485 33643
rect 15485 33609 15519 33643
rect 15519 33609 15528 33643
rect 15476 33600 15528 33609
rect 17960 33600 18012 33652
rect 22376 33643 22428 33652
rect 22376 33609 22385 33643
rect 22385 33609 22419 33643
rect 22419 33609 22428 33643
rect 22376 33600 22428 33609
rect 23572 33600 23624 33652
rect 24124 33600 24176 33652
rect 28632 33643 28684 33652
rect 28632 33609 28641 33643
rect 28641 33609 28675 33643
rect 28675 33609 28684 33643
rect 28632 33600 28684 33609
rect 30932 33600 30984 33652
rect 32588 33600 32640 33652
rect 33416 33643 33468 33652
rect 33416 33609 33425 33643
rect 33425 33609 33459 33643
rect 33459 33609 33468 33643
rect 33416 33600 33468 33609
rect 33508 33600 33560 33652
rect 2228 33464 2280 33516
rect 14372 33464 14424 33516
rect 17040 33532 17092 33584
rect 17868 33532 17920 33584
rect 21272 33532 21324 33584
rect 22284 33575 22336 33584
rect 22284 33541 22293 33575
rect 22293 33541 22327 33575
rect 22327 33541 22336 33575
rect 22284 33532 22336 33541
rect 25136 33532 25188 33584
rect 17500 33507 17552 33516
rect 17500 33473 17509 33507
rect 17509 33473 17543 33507
rect 17543 33473 17552 33507
rect 17500 33464 17552 33473
rect 17684 33507 17736 33516
rect 17684 33473 17693 33507
rect 17693 33473 17727 33507
rect 17727 33473 17736 33507
rect 17684 33464 17736 33473
rect 19340 33464 19392 33516
rect 23572 33464 23624 33516
rect 17132 33396 17184 33448
rect 22100 33396 22152 33448
rect 22468 33396 22520 33448
rect 23848 33507 23900 33516
rect 23848 33473 23857 33507
rect 23857 33473 23891 33507
rect 23891 33473 23900 33507
rect 23848 33464 23900 33473
rect 24032 33507 24084 33516
rect 24032 33473 24041 33507
rect 24041 33473 24075 33507
rect 24075 33473 24084 33507
rect 25412 33507 25464 33516
rect 24032 33464 24084 33473
rect 25412 33473 25421 33507
rect 25421 33473 25455 33507
rect 25455 33473 25464 33507
rect 25412 33464 25464 33473
rect 27160 33532 27212 33584
rect 24308 33396 24360 33448
rect 20444 33328 20496 33380
rect 23480 33328 23532 33380
rect 25044 33328 25096 33380
rect 28908 33464 28960 33516
rect 28356 33396 28408 33448
rect 29368 33464 29420 33516
rect 29552 33532 29604 33584
rect 31760 33532 31812 33584
rect 2872 33303 2924 33312
rect 2872 33269 2881 33303
rect 2881 33269 2915 33303
rect 2915 33269 2924 33303
rect 2872 33260 2924 33269
rect 17224 33260 17276 33312
rect 24032 33260 24084 33312
rect 25872 33260 25924 33312
rect 25964 33260 26016 33312
rect 27160 33260 27212 33312
rect 29828 33396 29880 33448
rect 30380 33507 30432 33516
rect 30380 33473 30414 33507
rect 30414 33473 30432 33507
rect 30380 33464 30432 33473
rect 40868 33532 40920 33584
rect 46480 33600 46532 33652
rect 31208 33328 31260 33380
rect 31484 33303 31536 33312
rect 31484 33269 31493 33303
rect 31493 33269 31527 33303
rect 31527 33269 31536 33303
rect 32588 33507 32640 33516
rect 32588 33473 32597 33507
rect 32597 33473 32631 33507
rect 32631 33473 32640 33507
rect 32772 33507 32824 33516
rect 32588 33464 32640 33473
rect 32772 33473 32781 33507
rect 32781 33473 32815 33507
rect 32815 33473 32824 33507
rect 32772 33464 32824 33473
rect 33324 33507 33376 33516
rect 33324 33473 33333 33507
rect 33333 33473 33367 33507
rect 33367 33473 33376 33507
rect 33324 33464 33376 33473
rect 45928 33507 45980 33516
rect 45928 33473 45937 33507
rect 45937 33473 45971 33507
rect 45971 33473 45980 33507
rect 45928 33464 45980 33473
rect 46572 33507 46624 33516
rect 46572 33473 46581 33507
rect 46581 33473 46615 33507
rect 46615 33473 46624 33507
rect 46572 33464 46624 33473
rect 47952 33507 48004 33516
rect 47952 33473 47961 33507
rect 47961 33473 47995 33507
rect 47995 33473 48004 33507
rect 47952 33464 48004 33473
rect 31484 33260 31536 33269
rect 46480 33260 46532 33312
rect 47952 33260 48004 33312
rect 48320 33260 48372 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 13268 32963 13320 32972
rect 13268 32929 13277 32963
rect 13277 32929 13311 32963
rect 13311 32929 13320 32963
rect 13268 32920 13320 32929
rect 1768 32852 1820 32904
rect 2596 32852 2648 32904
rect 3976 32852 4028 32904
rect 13912 32988 13964 33040
rect 13820 32852 13872 32904
rect 17684 32988 17736 33040
rect 15568 32920 15620 32972
rect 14740 32895 14792 32904
rect 14740 32861 14749 32895
rect 14749 32861 14783 32895
rect 14783 32861 14792 32895
rect 14740 32852 14792 32861
rect 16948 32852 17000 32904
rect 18144 32852 18196 32904
rect 19156 32852 19208 32904
rect 20812 32920 20864 32972
rect 16672 32827 16724 32836
rect 16672 32793 16706 32827
rect 16706 32793 16724 32827
rect 16672 32784 16724 32793
rect 19432 32784 19484 32836
rect 20444 32852 20496 32904
rect 21824 32920 21876 32972
rect 23572 33056 23624 33108
rect 24308 33056 24360 33108
rect 27160 33031 27212 33040
rect 27160 32997 27169 33031
rect 27169 32997 27203 33031
rect 27203 32997 27212 33031
rect 27160 32988 27212 32997
rect 29092 32988 29144 33040
rect 29368 32988 29420 33040
rect 32772 33056 32824 33108
rect 23572 32920 23624 32972
rect 24308 32920 24360 32972
rect 24676 32920 24728 32972
rect 29828 32920 29880 32972
rect 37004 32963 37056 32972
rect 37004 32929 37013 32963
rect 37013 32929 37047 32963
rect 37047 32929 37056 32963
rect 37004 32920 37056 32929
rect 46296 32963 46348 32972
rect 46296 32929 46305 32963
rect 46305 32929 46339 32963
rect 46339 32929 46348 32963
rect 46296 32920 46348 32929
rect 46480 32963 46532 32972
rect 46480 32929 46489 32963
rect 46489 32929 46523 32963
rect 46523 32929 46532 32963
rect 46480 32920 46532 32929
rect 48044 32963 48096 32972
rect 48044 32929 48053 32963
rect 48053 32929 48087 32963
rect 48087 32929 48096 32963
rect 48044 32920 48096 32929
rect 25780 32895 25832 32904
rect 20168 32784 20220 32836
rect 22008 32784 22060 32836
rect 22928 32784 22980 32836
rect 23296 32784 23348 32836
rect 1768 32716 1820 32768
rect 3056 32759 3108 32768
rect 3056 32725 3065 32759
rect 3065 32725 3099 32759
rect 3099 32725 3108 32759
rect 3056 32716 3108 32725
rect 14096 32759 14148 32768
rect 14096 32725 14105 32759
rect 14105 32725 14139 32759
rect 14139 32725 14148 32759
rect 14096 32716 14148 32725
rect 14464 32716 14516 32768
rect 19984 32716 20036 32768
rect 20720 32759 20772 32768
rect 20720 32725 20729 32759
rect 20729 32725 20763 32759
rect 20763 32725 20772 32759
rect 20720 32716 20772 32725
rect 21088 32759 21140 32768
rect 21088 32725 21097 32759
rect 21097 32725 21131 32759
rect 21131 32725 21140 32759
rect 21088 32716 21140 32725
rect 22192 32716 22244 32768
rect 23112 32716 23164 32768
rect 25780 32861 25789 32895
rect 25789 32861 25823 32895
rect 25823 32861 25832 32895
rect 25780 32852 25832 32861
rect 25872 32852 25924 32904
rect 26976 32852 27028 32904
rect 28540 32852 28592 32904
rect 27896 32827 27948 32836
rect 27896 32793 27905 32827
rect 27905 32793 27939 32827
rect 27939 32793 27948 32827
rect 27896 32784 27948 32793
rect 28908 32852 28960 32904
rect 29000 32895 29052 32904
rect 29000 32861 29009 32895
rect 29009 32861 29043 32895
rect 29043 32861 29052 32895
rect 29000 32852 29052 32861
rect 29736 32852 29788 32904
rect 31484 32852 31536 32904
rect 33876 32852 33928 32904
rect 29184 32784 29236 32836
rect 29460 32784 29512 32836
rect 30288 32784 30340 32836
rect 32404 32827 32456 32836
rect 32404 32793 32413 32827
rect 32413 32793 32447 32827
rect 32447 32793 32456 32827
rect 32404 32784 32456 32793
rect 35348 32827 35400 32836
rect 35348 32793 35357 32827
rect 35357 32793 35391 32827
rect 35391 32793 35400 32827
rect 35348 32784 35400 32793
rect 25964 32716 26016 32768
rect 30012 32759 30064 32768
rect 30012 32725 30021 32759
rect 30021 32725 30055 32759
rect 30055 32725 30064 32759
rect 30012 32716 30064 32725
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 10968 32512 11020 32564
rect 13268 32512 13320 32564
rect 16672 32555 16724 32564
rect 16672 32521 16681 32555
rect 16681 32521 16715 32555
rect 16715 32521 16724 32555
rect 16672 32512 16724 32521
rect 17868 32512 17920 32564
rect 21088 32512 21140 32564
rect 24952 32512 25004 32564
rect 25320 32555 25372 32564
rect 25320 32521 25329 32555
rect 25329 32521 25363 32555
rect 25363 32521 25372 32555
rect 25320 32512 25372 32521
rect 26332 32555 26384 32564
rect 26332 32521 26341 32555
rect 26341 32521 26375 32555
rect 26375 32521 26384 32555
rect 26332 32512 26384 32521
rect 14096 32444 14148 32496
rect 1768 32419 1820 32428
rect 1768 32385 1777 32419
rect 1777 32385 1811 32419
rect 1811 32385 1820 32419
rect 1768 32376 1820 32385
rect 10876 32376 10928 32428
rect 1952 32351 2004 32360
rect 1952 32317 1961 32351
rect 1961 32317 1995 32351
rect 1995 32317 2004 32351
rect 1952 32308 2004 32317
rect 2780 32351 2832 32360
rect 2780 32317 2789 32351
rect 2789 32317 2823 32351
rect 2823 32317 2832 32351
rect 2780 32308 2832 32317
rect 14280 32376 14332 32428
rect 16580 32376 16632 32428
rect 14004 32308 14056 32360
rect 17224 32376 17276 32428
rect 17592 32444 17644 32496
rect 18144 32487 18196 32496
rect 18144 32453 18153 32487
rect 18153 32453 18187 32487
rect 18187 32453 18196 32487
rect 18144 32444 18196 32453
rect 17868 32419 17920 32428
rect 17868 32385 17877 32419
rect 17877 32385 17911 32419
rect 17911 32385 17920 32419
rect 17868 32376 17920 32385
rect 18052 32419 18104 32428
rect 18052 32385 18061 32419
rect 18061 32385 18095 32419
rect 18095 32385 18104 32419
rect 18052 32376 18104 32385
rect 20628 32444 20680 32496
rect 19892 32419 19944 32428
rect 19892 32385 19926 32419
rect 19926 32385 19944 32419
rect 19892 32376 19944 32385
rect 22284 32444 22336 32496
rect 23848 32444 23900 32496
rect 21916 32376 21968 32428
rect 24032 32376 24084 32428
rect 25780 32444 25832 32496
rect 25688 32376 25740 32428
rect 24952 32308 25004 32360
rect 26240 32376 26292 32428
rect 12716 32172 12768 32224
rect 17132 32240 17184 32292
rect 27344 32308 27396 32360
rect 30012 32512 30064 32564
rect 27896 32444 27948 32496
rect 33876 32444 33928 32496
rect 28448 32376 28500 32428
rect 28632 32376 28684 32428
rect 29000 32376 29052 32428
rect 31852 32376 31904 32428
rect 32404 32419 32456 32428
rect 32404 32385 32413 32419
rect 32413 32385 32447 32419
rect 32447 32385 32456 32419
rect 32404 32376 32456 32385
rect 29644 32351 29696 32360
rect 13912 32172 13964 32224
rect 22928 32172 22980 32224
rect 28908 32240 28960 32292
rect 29644 32317 29653 32351
rect 29653 32317 29687 32351
rect 29687 32317 29696 32351
rect 29644 32308 29696 32317
rect 29828 32351 29880 32360
rect 29828 32317 29837 32351
rect 29837 32317 29871 32351
rect 29871 32317 29880 32351
rect 29828 32308 29880 32317
rect 30104 32308 30156 32360
rect 31760 32240 31812 32292
rect 25320 32172 25372 32224
rect 26148 32172 26200 32224
rect 26792 32172 26844 32224
rect 28632 32172 28684 32224
rect 30196 32172 30248 32224
rect 32772 32172 32824 32224
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4068 31968 4120 32020
rect 10876 32011 10928 32020
rect 2964 31900 3016 31952
rect 10876 31977 10885 32011
rect 10885 31977 10919 32011
rect 10919 31977 10928 32011
rect 10876 31968 10928 31977
rect 21916 32011 21968 32020
rect 11244 31900 11296 31952
rect 13176 31900 13228 31952
rect 21916 31977 21925 32011
rect 21925 31977 21959 32011
rect 21959 31977 21968 32011
rect 21916 31968 21968 31977
rect 25688 31968 25740 32020
rect 10140 31875 10192 31884
rect 10140 31841 10149 31875
rect 10149 31841 10183 31875
rect 10183 31841 10192 31875
rect 10140 31832 10192 31841
rect 3240 31807 3292 31816
rect 3240 31773 3249 31807
rect 3249 31773 3283 31807
rect 3283 31773 3292 31807
rect 3240 31764 3292 31773
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 10876 31764 10928 31816
rect 11152 31807 11204 31816
rect 11152 31773 11161 31807
rect 11161 31773 11195 31807
rect 11195 31773 11204 31807
rect 11152 31764 11204 31773
rect 14372 31875 14424 31884
rect 14372 31841 14381 31875
rect 14381 31841 14415 31875
rect 14415 31841 14424 31875
rect 14372 31832 14424 31841
rect 11520 31807 11572 31816
rect 11520 31773 11529 31807
rect 11529 31773 11563 31807
rect 11563 31773 11572 31807
rect 11520 31764 11572 31773
rect 12716 31764 12768 31816
rect 17960 31832 18012 31884
rect 19340 31832 19392 31884
rect 20260 31832 20312 31884
rect 21088 31832 21140 31884
rect 17224 31807 17276 31816
rect 17224 31773 17233 31807
rect 17233 31773 17267 31807
rect 17267 31773 17276 31807
rect 17224 31764 17276 31773
rect 17868 31807 17920 31816
rect 13084 31696 13136 31748
rect 17868 31773 17877 31807
rect 17877 31773 17911 31807
rect 17911 31773 17920 31807
rect 17868 31764 17920 31773
rect 20996 31764 21048 31816
rect 22652 31832 22704 31884
rect 26332 31832 26384 31884
rect 22376 31801 22428 31816
rect 22376 31767 22408 31801
rect 22408 31767 22428 31801
rect 22376 31764 22428 31767
rect 23480 31764 23532 31816
rect 25228 31764 25280 31816
rect 26240 31764 26292 31816
rect 27160 31832 27212 31884
rect 28356 31968 28408 32020
rect 29736 31968 29788 32020
rect 31852 31968 31904 32020
rect 33876 32011 33928 32020
rect 33876 31977 33885 32011
rect 33885 31977 33919 32011
rect 33919 31977 33928 32011
rect 33876 31968 33928 31977
rect 34336 31968 34388 32020
rect 35348 32011 35400 32020
rect 35348 31977 35357 32011
rect 35357 31977 35391 32011
rect 35391 31977 35400 32011
rect 35348 31968 35400 31977
rect 17960 31696 18012 31748
rect 19432 31696 19484 31748
rect 22008 31696 22060 31748
rect 25136 31696 25188 31748
rect 26792 31807 26844 31816
rect 26792 31773 26801 31807
rect 26801 31773 26835 31807
rect 26835 31773 26844 31807
rect 28908 31832 28960 31884
rect 29828 31832 29880 31884
rect 47860 31875 47912 31884
rect 47860 31841 47869 31875
rect 47869 31841 47903 31875
rect 47903 31841 47912 31875
rect 47860 31832 47912 31841
rect 26792 31764 26844 31773
rect 31760 31764 31812 31816
rect 37280 31764 37332 31816
rect 47492 31807 47544 31816
rect 47492 31773 47501 31807
rect 47501 31773 47535 31807
rect 47535 31773 47544 31807
rect 47492 31764 47544 31773
rect 14740 31628 14792 31680
rect 22468 31628 22520 31680
rect 25780 31628 25832 31680
rect 27160 31628 27212 31680
rect 28356 31696 28408 31748
rect 29552 31739 29604 31748
rect 29552 31705 29561 31739
rect 29561 31705 29595 31739
rect 29595 31705 29604 31739
rect 29552 31696 29604 31705
rect 29736 31739 29788 31748
rect 29736 31705 29745 31739
rect 29745 31705 29779 31739
rect 29779 31705 29788 31739
rect 29736 31696 29788 31705
rect 30472 31696 30524 31748
rect 32128 31696 32180 31748
rect 29092 31628 29144 31680
rect 30012 31628 30064 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 13084 31467 13136 31476
rect 13084 31433 13093 31467
rect 13093 31433 13127 31467
rect 13127 31433 13136 31467
rect 13084 31424 13136 31433
rect 13268 31424 13320 31476
rect 1492 31399 1544 31408
rect 1492 31365 1501 31399
rect 1501 31365 1535 31399
rect 1535 31365 1544 31399
rect 1492 31356 1544 31365
rect 3056 31356 3108 31408
rect 5264 31356 5316 31408
rect 12992 31356 13044 31408
rect 14096 31424 14148 31476
rect 14740 31356 14792 31408
rect 20260 31356 20312 31408
rect 20628 31356 20680 31408
rect 20996 31424 21048 31476
rect 13360 31331 13412 31340
rect 13360 31297 13369 31331
rect 13369 31297 13403 31331
rect 13403 31297 13412 31331
rect 13360 31288 13412 31297
rect 3148 31263 3200 31272
rect 3148 31229 3157 31263
rect 3157 31229 3191 31263
rect 3191 31229 3200 31263
rect 3148 31220 3200 31229
rect 13820 31263 13872 31272
rect 2872 31152 2924 31204
rect 13820 31229 13829 31263
rect 13829 31229 13863 31263
rect 13863 31229 13872 31263
rect 13820 31220 13872 31229
rect 14004 31288 14056 31340
rect 14372 31288 14424 31340
rect 16764 31288 16816 31340
rect 18788 31288 18840 31340
rect 19248 31288 19300 31340
rect 20996 31288 21048 31340
rect 15108 31220 15160 31272
rect 15200 31220 15252 31272
rect 20812 31220 20864 31272
rect 22376 31424 22428 31476
rect 22468 31424 22520 31476
rect 24308 31467 24360 31476
rect 22192 31356 22244 31408
rect 23296 31356 23348 31408
rect 24308 31433 24317 31467
rect 24317 31433 24351 31467
rect 24351 31433 24360 31467
rect 24308 31424 24360 31433
rect 26792 31424 26844 31476
rect 29552 31424 29604 31476
rect 30472 31424 30524 31476
rect 32128 31467 32180 31476
rect 32128 31433 32137 31467
rect 32137 31433 32171 31467
rect 32171 31433 32180 31467
rect 32128 31424 32180 31433
rect 24768 31356 24820 31408
rect 26240 31356 26292 31408
rect 26424 31356 26476 31408
rect 27896 31356 27948 31408
rect 28816 31356 28868 31408
rect 23020 31331 23072 31340
rect 23020 31297 23029 31331
rect 23029 31297 23063 31331
rect 23063 31297 23072 31331
rect 23020 31288 23072 31297
rect 24032 31288 24084 31340
rect 24400 31288 24452 31340
rect 23112 31220 23164 31272
rect 23848 31220 23900 31272
rect 25044 31220 25096 31272
rect 12716 31152 12768 31204
rect 20168 31152 20220 31204
rect 21364 31152 21416 31204
rect 29644 31288 29696 31340
rect 26148 31220 26200 31272
rect 13728 31127 13780 31136
rect 13728 31093 13737 31127
rect 13737 31093 13771 31127
rect 13771 31093 13780 31127
rect 13728 31084 13780 31093
rect 14464 31084 14516 31136
rect 18052 31127 18104 31136
rect 18052 31093 18061 31127
rect 18061 31093 18095 31127
rect 18095 31093 18104 31127
rect 18052 31084 18104 31093
rect 19248 31084 19300 31136
rect 23296 31084 23348 31136
rect 25964 31127 26016 31136
rect 25964 31093 25973 31127
rect 25973 31093 26007 31127
rect 26007 31093 26016 31127
rect 25964 31084 26016 31093
rect 26976 31084 27028 31136
rect 27160 31127 27212 31136
rect 27160 31093 27169 31127
rect 27169 31093 27203 31127
rect 27203 31093 27212 31127
rect 27160 31084 27212 31093
rect 28908 31152 28960 31204
rect 29736 31220 29788 31272
rect 30196 31331 30248 31340
rect 30196 31297 30205 31331
rect 30205 31297 30239 31331
rect 30239 31297 30248 31331
rect 30196 31288 30248 31297
rect 30380 31331 30432 31340
rect 30380 31297 30389 31331
rect 30389 31297 30423 31331
rect 30423 31297 30432 31331
rect 30380 31288 30432 31297
rect 31852 31356 31904 31408
rect 30932 31288 30984 31340
rect 32588 31331 32640 31340
rect 32588 31297 32597 31331
rect 32597 31297 32631 31331
rect 32631 31297 32640 31331
rect 32772 31331 32824 31340
rect 32588 31288 32640 31297
rect 32772 31297 32781 31331
rect 32781 31297 32815 31331
rect 32815 31297 32824 31331
rect 32772 31288 32824 31297
rect 47952 31331 48004 31340
rect 47952 31297 47961 31331
rect 47961 31297 47995 31331
rect 47995 31297 48004 31331
rect 47952 31288 48004 31297
rect 30196 31152 30248 31204
rect 38844 31152 38896 31204
rect 29184 31084 29236 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 1952 30880 2004 30932
rect 2964 30880 3016 30932
rect 10140 30880 10192 30932
rect 16856 30923 16908 30932
rect 16856 30889 16865 30923
rect 16865 30889 16899 30923
rect 16899 30889 16908 30923
rect 16856 30880 16908 30889
rect 17868 30880 17920 30932
rect 23020 30880 23072 30932
rect 24768 30880 24820 30932
rect 11244 30812 11296 30864
rect 11796 30812 11848 30864
rect 15200 30855 15252 30864
rect 15200 30821 15209 30855
rect 15209 30821 15243 30855
rect 15243 30821 15252 30855
rect 15200 30812 15252 30821
rect 20444 30812 20496 30864
rect 2964 30676 3016 30728
rect 10048 30676 10100 30728
rect 10416 30719 10468 30728
rect 10416 30685 10425 30719
rect 10425 30685 10459 30719
rect 10459 30685 10468 30719
rect 10416 30676 10468 30685
rect 11152 30719 11204 30728
rect 11152 30685 11161 30719
rect 11161 30685 11195 30719
rect 11195 30685 11204 30719
rect 11152 30676 11204 30685
rect 11520 30719 11572 30728
rect 8300 30608 8352 30660
rect 9956 30540 10008 30592
rect 11520 30685 11529 30719
rect 11529 30685 11563 30719
rect 11563 30685 11572 30719
rect 11520 30676 11572 30685
rect 13912 30676 13964 30728
rect 14280 30719 14332 30728
rect 14280 30685 14289 30719
rect 14289 30685 14323 30719
rect 14323 30685 14332 30719
rect 14280 30676 14332 30685
rect 17408 30676 17460 30728
rect 18052 30744 18104 30796
rect 20168 30744 20220 30796
rect 23480 30812 23532 30864
rect 24308 30812 24360 30864
rect 21824 30744 21876 30796
rect 24860 30787 24912 30796
rect 24860 30753 24869 30787
rect 24869 30753 24903 30787
rect 24903 30753 24912 30787
rect 24860 30744 24912 30753
rect 25504 30812 25556 30864
rect 25872 30812 25924 30864
rect 25964 30812 26016 30864
rect 17224 30608 17276 30660
rect 20168 30608 20220 30660
rect 22100 30676 22152 30728
rect 23112 30719 23164 30728
rect 23112 30685 23121 30719
rect 23121 30685 23155 30719
rect 23155 30685 23164 30719
rect 23112 30676 23164 30685
rect 21272 30608 21324 30660
rect 21364 30608 21416 30660
rect 23296 30719 23348 30728
rect 23296 30685 23305 30719
rect 23305 30685 23339 30719
rect 23339 30685 23348 30719
rect 23296 30676 23348 30685
rect 23480 30719 23532 30728
rect 23480 30685 23489 30719
rect 23489 30685 23523 30719
rect 23523 30685 23532 30719
rect 23480 30676 23532 30685
rect 25780 30676 25832 30728
rect 26056 30719 26108 30728
rect 26056 30685 26065 30719
rect 26065 30685 26099 30719
rect 26099 30685 26108 30719
rect 26792 30880 26844 30932
rect 30196 30880 30248 30932
rect 41512 30880 41564 30932
rect 26056 30676 26108 30685
rect 26332 30676 26384 30728
rect 26976 30719 27028 30728
rect 26976 30685 26985 30719
rect 26985 30685 27019 30719
rect 27019 30685 27028 30719
rect 26976 30676 27028 30685
rect 29184 30676 29236 30728
rect 42800 30744 42852 30796
rect 25136 30608 25188 30660
rect 26424 30608 26476 30660
rect 30012 30719 30064 30728
rect 30012 30685 30021 30719
rect 30021 30685 30055 30719
rect 30055 30685 30064 30719
rect 30012 30676 30064 30685
rect 30288 30676 30340 30728
rect 33232 30719 33284 30728
rect 33232 30685 33241 30719
rect 33241 30685 33275 30719
rect 33275 30685 33284 30719
rect 33232 30676 33284 30685
rect 33508 30676 33560 30728
rect 33968 30719 34020 30728
rect 33968 30685 33977 30719
rect 33977 30685 34011 30719
rect 34011 30685 34020 30719
rect 33968 30676 34020 30685
rect 34336 30676 34388 30728
rect 40132 30676 40184 30728
rect 14372 30540 14424 30592
rect 16948 30540 17000 30592
rect 17684 30583 17736 30592
rect 17684 30549 17693 30583
rect 17693 30549 17727 30583
rect 17727 30549 17736 30583
rect 17684 30540 17736 30549
rect 19432 30583 19484 30592
rect 19432 30549 19441 30583
rect 19441 30549 19475 30583
rect 19475 30549 19484 30583
rect 19432 30540 19484 30549
rect 20812 30540 20864 30592
rect 21640 30583 21692 30592
rect 21640 30549 21649 30583
rect 21649 30549 21683 30583
rect 21683 30549 21692 30583
rect 21640 30540 21692 30549
rect 22744 30540 22796 30592
rect 23020 30540 23072 30592
rect 24308 30540 24360 30592
rect 25596 30583 25648 30592
rect 25596 30549 25605 30583
rect 25605 30549 25639 30583
rect 25639 30549 25648 30583
rect 25596 30540 25648 30549
rect 29092 30540 29144 30592
rect 29184 30540 29236 30592
rect 33416 30608 33468 30660
rect 48504 30608 48556 30660
rect 31668 30540 31720 30592
rect 32220 30540 32272 30592
rect 33600 30540 33652 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 9680 30336 9732 30388
rect 10416 30336 10468 30388
rect 10968 30379 11020 30388
rect 10968 30345 10977 30379
rect 10977 30345 11011 30379
rect 11011 30345 11020 30379
rect 10968 30336 11020 30345
rect 13360 30336 13412 30388
rect 18512 30336 18564 30388
rect 21272 30379 21324 30388
rect 21272 30345 21281 30379
rect 21281 30345 21315 30379
rect 21315 30345 21324 30379
rect 21272 30336 21324 30345
rect 23480 30336 23532 30388
rect 24952 30379 25004 30388
rect 24952 30345 24961 30379
rect 24961 30345 24995 30379
rect 24995 30345 25004 30379
rect 24952 30336 25004 30345
rect 26056 30336 26108 30388
rect 29092 30336 29144 30388
rect 2044 30200 2096 30252
rect 8208 30268 8260 30320
rect 8300 30200 8352 30252
rect 12716 30268 12768 30320
rect 10324 30200 10376 30252
rect 11152 30200 11204 30252
rect 14372 30268 14424 30320
rect 17040 30268 17092 30320
rect 21640 30268 21692 30320
rect 11428 30132 11480 30184
rect 14464 30243 14516 30252
rect 13820 30175 13872 30184
rect 13820 30141 13829 30175
rect 13829 30141 13863 30175
rect 13863 30141 13872 30175
rect 13820 30132 13872 30141
rect 13728 30107 13780 30116
rect 13728 30073 13737 30107
rect 13737 30073 13771 30107
rect 13771 30073 13780 30107
rect 13728 30064 13780 30073
rect 14464 30209 14473 30243
rect 14473 30209 14507 30243
rect 14507 30209 14516 30243
rect 14464 30200 14516 30209
rect 14004 30132 14056 30184
rect 1400 29996 1452 30048
rect 2320 30039 2372 30048
rect 2320 30005 2329 30039
rect 2329 30005 2363 30039
rect 2363 30005 2372 30039
rect 2320 29996 2372 30005
rect 9312 29996 9364 30048
rect 13084 30039 13136 30048
rect 13084 30005 13093 30039
rect 13093 30005 13127 30039
rect 13127 30005 13136 30039
rect 13084 29996 13136 30005
rect 14464 29996 14516 30048
rect 16580 30200 16632 30252
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 17500 30243 17552 30252
rect 16948 30200 17000 30209
rect 17500 30209 17509 30243
rect 17509 30209 17543 30243
rect 17543 30209 17552 30243
rect 17500 30200 17552 30209
rect 19432 30200 19484 30252
rect 20996 30200 21048 30252
rect 26332 30268 26384 30320
rect 31392 30336 31444 30388
rect 23020 30200 23072 30252
rect 23572 30200 23624 30252
rect 17408 30132 17460 30184
rect 18420 30175 18472 30184
rect 18420 30141 18429 30175
rect 18429 30141 18463 30175
rect 18463 30141 18472 30175
rect 18420 30132 18472 30141
rect 25044 30200 25096 30252
rect 25412 30200 25464 30252
rect 30932 30200 30984 30252
rect 33600 30311 33652 30320
rect 33600 30277 33609 30311
rect 33609 30277 33643 30311
rect 33643 30277 33652 30311
rect 33600 30268 33652 30277
rect 25780 30132 25832 30184
rect 29276 30132 29328 30184
rect 31668 30200 31720 30252
rect 31944 30200 31996 30252
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 33232 30200 33284 30252
rect 35440 30132 35492 30184
rect 16580 30064 16632 30116
rect 16764 30064 16816 30116
rect 18052 29996 18104 30048
rect 18144 29996 18196 30048
rect 22744 29996 22796 30048
rect 24308 30039 24360 30048
rect 24308 30005 24317 30039
rect 24317 30005 24351 30039
rect 24351 30005 24360 30039
rect 24308 29996 24360 30005
rect 25044 29996 25096 30048
rect 35532 30064 35584 30116
rect 31852 29996 31904 30048
rect 31944 29996 31996 30048
rect 32312 29996 32364 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 10324 29835 10376 29844
rect 10324 29801 10333 29835
rect 10333 29801 10367 29835
rect 10367 29801 10376 29835
rect 10324 29792 10376 29801
rect 10968 29792 11020 29844
rect 6368 29724 6420 29776
rect 1400 29699 1452 29708
rect 1400 29665 1409 29699
rect 1409 29665 1443 29699
rect 1443 29665 1452 29699
rect 1400 29656 1452 29665
rect 2320 29656 2372 29708
rect 2780 29699 2832 29708
rect 2780 29665 2789 29699
rect 2789 29665 2823 29699
rect 2823 29665 2832 29699
rect 2780 29656 2832 29665
rect 11796 29699 11848 29708
rect 10048 29588 10100 29640
rect 10600 29631 10652 29640
rect 10600 29597 10609 29631
rect 10609 29597 10643 29631
rect 10643 29597 10652 29631
rect 10600 29588 10652 29597
rect 11796 29665 11805 29699
rect 11805 29665 11839 29699
rect 11839 29665 11848 29699
rect 11796 29656 11848 29665
rect 13728 29656 13780 29708
rect 13912 29656 13964 29708
rect 9680 29563 9732 29572
rect 9680 29529 9689 29563
rect 9689 29529 9723 29563
rect 9723 29529 9732 29563
rect 9680 29520 9732 29529
rect 11336 29588 11388 29640
rect 11428 29520 11480 29572
rect 10140 29452 10192 29504
rect 10876 29452 10928 29504
rect 17684 29724 17736 29776
rect 17408 29588 17460 29640
rect 18144 29792 18196 29844
rect 18420 29792 18472 29844
rect 18512 29792 18564 29844
rect 23756 29792 23808 29844
rect 25412 29792 25464 29844
rect 32128 29792 32180 29844
rect 34520 29792 34572 29844
rect 22744 29724 22796 29776
rect 25780 29724 25832 29776
rect 31668 29724 31720 29776
rect 19248 29656 19300 29708
rect 27344 29656 27396 29708
rect 28172 29699 28224 29708
rect 28172 29665 28181 29699
rect 28181 29665 28215 29699
rect 28215 29665 28224 29699
rect 28172 29656 28224 29665
rect 28448 29656 28500 29708
rect 14280 29520 14332 29572
rect 15844 29563 15896 29572
rect 15844 29529 15853 29563
rect 15853 29529 15887 29563
rect 15887 29529 15896 29563
rect 15844 29520 15896 29529
rect 16028 29563 16080 29572
rect 16028 29529 16037 29563
rect 16037 29529 16071 29563
rect 16071 29529 16080 29563
rect 16028 29520 16080 29529
rect 15292 29495 15344 29504
rect 15292 29461 15301 29495
rect 15301 29461 15335 29495
rect 15335 29461 15344 29495
rect 15292 29452 15344 29461
rect 15936 29452 15988 29504
rect 16304 29452 16356 29504
rect 18052 29631 18104 29640
rect 18052 29597 18061 29631
rect 18061 29597 18095 29631
rect 18095 29597 18104 29631
rect 18052 29588 18104 29597
rect 19432 29588 19484 29640
rect 20812 29588 20864 29640
rect 26332 29588 26384 29640
rect 27252 29588 27304 29640
rect 27804 29588 27856 29640
rect 30932 29631 30984 29640
rect 30932 29597 30941 29631
rect 30941 29597 30975 29631
rect 30975 29597 30984 29631
rect 30932 29588 30984 29597
rect 31208 29656 31260 29708
rect 31760 29699 31812 29708
rect 31760 29665 31769 29699
rect 31769 29665 31803 29699
rect 31803 29665 31812 29699
rect 35532 29699 35584 29708
rect 31760 29656 31812 29665
rect 35532 29665 35541 29699
rect 35541 29665 35575 29699
rect 35575 29665 35584 29699
rect 35532 29656 35584 29665
rect 42800 29656 42852 29708
rect 19340 29520 19392 29572
rect 20628 29520 20680 29572
rect 25596 29520 25648 29572
rect 18696 29452 18748 29504
rect 22192 29452 22244 29504
rect 24308 29452 24360 29504
rect 31392 29520 31444 29572
rect 31852 29588 31904 29640
rect 33508 29588 33560 29640
rect 33968 29588 34020 29640
rect 34612 29588 34664 29640
rect 47308 29631 47360 29640
rect 47308 29597 47317 29631
rect 47317 29597 47351 29631
rect 47351 29597 47360 29631
rect 47308 29588 47360 29597
rect 32220 29520 32272 29572
rect 35716 29563 35768 29572
rect 35716 29529 35725 29563
rect 35725 29529 35759 29563
rect 35759 29529 35768 29563
rect 35716 29520 35768 29529
rect 46848 29520 46900 29572
rect 27712 29452 27764 29504
rect 32128 29452 32180 29504
rect 33692 29495 33744 29504
rect 33692 29461 33701 29495
rect 33701 29461 33735 29495
rect 33735 29461 33744 29495
rect 33692 29452 33744 29461
rect 34796 29495 34848 29504
rect 34796 29461 34805 29495
rect 34805 29461 34839 29495
rect 34839 29461 34848 29495
rect 34796 29452 34848 29461
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 9956 29291 10008 29300
rect 9956 29257 9965 29291
rect 9965 29257 9999 29291
rect 9999 29257 10008 29291
rect 9956 29248 10008 29257
rect 10048 29248 10100 29300
rect 11796 29248 11848 29300
rect 14464 29248 14516 29300
rect 15292 29248 15344 29300
rect 9220 29180 9272 29232
rect 2688 29112 2740 29164
rect 2964 29155 3016 29164
rect 2964 29121 2973 29155
rect 2973 29121 3007 29155
rect 3007 29121 3016 29155
rect 2964 29112 3016 29121
rect 10048 29155 10100 29164
rect 10048 29121 10057 29155
rect 10057 29121 10091 29155
rect 10091 29121 10100 29155
rect 10048 29112 10100 29121
rect 13084 29180 13136 29232
rect 12716 29155 12768 29164
rect 12716 29121 12725 29155
rect 12725 29121 12759 29155
rect 12759 29121 12768 29155
rect 12716 29112 12768 29121
rect 16488 29180 16540 29232
rect 12624 29044 12676 29096
rect 14096 29019 14148 29028
rect 14096 28985 14105 29019
rect 14105 28985 14139 29019
rect 14139 28985 14148 29019
rect 15660 29044 15712 29096
rect 15936 29155 15988 29164
rect 15936 29121 15945 29155
rect 15945 29121 15979 29155
rect 15979 29121 15988 29155
rect 15936 29112 15988 29121
rect 16120 29155 16172 29164
rect 16120 29121 16129 29155
rect 16129 29121 16163 29155
rect 16163 29121 16172 29155
rect 16120 29112 16172 29121
rect 16304 29112 16356 29164
rect 19432 29180 19484 29232
rect 17316 29112 17368 29164
rect 17868 29112 17920 29164
rect 21088 29112 21140 29164
rect 22192 29248 22244 29300
rect 23572 29223 23624 29232
rect 23572 29189 23581 29223
rect 23581 29189 23615 29223
rect 23615 29189 23624 29223
rect 23572 29180 23624 29189
rect 23756 29180 23808 29232
rect 28448 29180 28500 29232
rect 29000 29180 29052 29232
rect 14096 28976 14148 28985
rect 1860 28951 1912 28960
rect 1860 28917 1869 28951
rect 1869 28917 1903 28951
rect 1903 28917 1912 28951
rect 1860 28908 1912 28917
rect 2412 28951 2464 28960
rect 2412 28917 2421 28951
rect 2421 28917 2455 28951
rect 2455 28917 2464 28951
rect 2412 28908 2464 28917
rect 2872 28908 2924 28960
rect 11244 28908 11296 28960
rect 23112 29044 23164 29096
rect 29184 29112 29236 29164
rect 29644 29248 29696 29300
rect 29828 29248 29880 29300
rect 33416 29248 33468 29300
rect 35716 29248 35768 29300
rect 29368 29180 29420 29232
rect 32128 29180 32180 29232
rect 31392 29112 31444 29164
rect 25780 29087 25832 29096
rect 18052 29019 18104 29028
rect 18052 28985 18061 29019
rect 18061 28985 18095 29019
rect 18095 28985 18104 29019
rect 18052 28976 18104 28985
rect 25044 28976 25096 29028
rect 25780 29053 25789 29087
rect 25789 29053 25823 29087
rect 25823 29053 25832 29087
rect 25780 29044 25832 29053
rect 31760 29112 31812 29164
rect 37464 29180 37516 29232
rect 34520 29155 34572 29164
rect 32128 29044 32180 29096
rect 34520 29121 34529 29155
rect 34529 29121 34563 29155
rect 34563 29121 34572 29155
rect 34520 29112 34572 29121
rect 37280 29155 37332 29164
rect 37280 29121 37289 29155
rect 37289 29121 37323 29155
rect 37323 29121 37332 29155
rect 37280 29112 37332 29121
rect 45836 29112 45888 29164
rect 47216 29112 47268 29164
rect 34704 29087 34756 29096
rect 34704 29053 34713 29087
rect 34713 29053 34747 29087
rect 34747 29053 34756 29087
rect 34704 29044 34756 29053
rect 36360 29087 36412 29096
rect 36360 29053 36369 29087
rect 36369 29053 36403 29087
rect 36403 29053 36412 29087
rect 36360 29044 36412 29053
rect 16580 28908 16632 28960
rect 17316 28908 17368 28960
rect 19340 28908 19392 28960
rect 23296 28908 23348 28960
rect 25872 28908 25924 28960
rect 34888 28976 34940 29028
rect 30840 28951 30892 28960
rect 30840 28917 30849 28951
rect 30849 28917 30883 28951
rect 30883 28917 30892 28951
rect 30840 28908 30892 28917
rect 34060 28908 34112 28960
rect 47032 28951 47084 28960
rect 47032 28917 47041 28951
rect 47041 28917 47075 28951
rect 47075 28917 47084 28951
rect 47032 28908 47084 28917
rect 47676 28951 47728 28960
rect 47676 28917 47685 28951
rect 47685 28917 47719 28951
rect 47719 28917 47728 28951
rect 47676 28908 47728 28917
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 1860 28568 1912 28620
rect 2780 28611 2832 28620
rect 2780 28577 2789 28611
rect 2789 28577 2823 28611
rect 2823 28577 2832 28611
rect 2780 28568 2832 28577
rect 9128 28500 9180 28552
rect 10048 28704 10100 28756
rect 10876 28704 10928 28756
rect 17316 28747 17368 28756
rect 17316 28713 17325 28747
rect 17325 28713 17359 28747
rect 17359 28713 17368 28747
rect 17316 28704 17368 28713
rect 17408 28704 17460 28756
rect 9496 28636 9548 28688
rect 11152 28636 11204 28688
rect 11336 28636 11388 28688
rect 11520 28636 11572 28688
rect 14740 28636 14792 28688
rect 18236 28704 18288 28756
rect 20076 28704 20128 28756
rect 20996 28704 21048 28756
rect 23756 28747 23808 28756
rect 23756 28713 23765 28747
rect 23765 28713 23799 28747
rect 23799 28713 23808 28747
rect 23756 28704 23808 28713
rect 24768 28704 24820 28756
rect 25504 28747 25556 28756
rect 25504 28713 25513 28747
rect 25513 28713 25547 28747
rect 25547 28713 25556 28747
rect 25504 28704 25556 28713
rect 27068 28704 27120 28756
rect 33232 28704 33284 28756
rect 34704 28704 34756 28756
rect 14004 28568 14056 28620
rect 14280 28611 14332 28620
rect 14280 28577 14289 28611
rect 14289 28577 14323 28611
rect 14323 28577 14332 28611
rect 14280 28568 14332 28577
rect 14464 28611 14516 28620
rect 14464 28577 14473 28611
rect 14473 28577 14507 28611
rect 14507 28577 14516 28611
rect 14464 28568 14516 28577
rect 9404 28543 9456 28552
rect 9404 28509 9413 28543
rect 9413 28509 9447 28543
rect 9447 28509 9456 28543
rect 9404 28500 9456 28509
rect 9588 28543 9640 28552
rect 9588 28509 9597 28543
rect 9597 28509 9631 28543
rect 9631 28509 9640 28543
rect 9588 28500 9640 28509
rect 10600 28500 10652 28552
rect 2412 28432 2464 28484
rect 8024 28475 8076 28484
rect 8024 28441 8033 28475
rect 8033 28441 8067 28475
rect 8067 28441 8076 28475
rect 8024 28432 8076 28441
rect 8576 28432 8628 28484
rect 11152 28432 11204 28484
rect 11336 28543 11388 28552
rect 11336 28509 11345 28543
rect 11345 28509 11379 28543
rect 11379 28509 11388 28543
rect 12072 28543 12124 28552
rect 11336 28500 11388 28509
rect 12072 28509 12081 28543
rect 12081 28509 12115 28543
rect 12115 28509 12124 28543
rect 12072 28500 12124 28509
rect 12440 28543 12492 28552
rect 12440 28509 12449 28543
rect 12449 28509 12483 28543
rect 12483 28509 12492 28543
rect 12440 28500 12492 28509
rect 12624 28500 12676 28552
rect 14372 28543 14424 28552
rect 14372 28509 14381 28543
rect 14381 28509 14415 28543
rect 14415 28509 14424 28543
rect 14372 28500 14424 28509
rect 14740 28500 14792 28552
rect 15844 28568 15896 28620
rect 16580 28568 16632 28620
rect 18052 28679 18104 28688
rect 18052 28645 18061 28679
rect 18061 28645 18095 28679
rect 18095 28645 18104 28679
rect 18052 28636 18104 28645
rect 25872 28636 25924 28688
rect 17592 28568 17644 28620
rect 19432 28611 19484 28620
rect 16488 28500 16540 28552
rect 18144 28500 18196 28552
rect 8484 28364 8536 28416
rect 10600 28407 10652 28416
rect 10600 28373 10609 28407
rect 10609 28373 10643 28407
rect 10643 28373 10652 28407
rect 10600 28364 10652 28373
rect 11060 28407 11112 28416
rect 11060 28373 11069 28407
rect 11069 28373 11103 28407
rect 11103 28373 11112 28407
rect 11060 28364 11112 28373
rect 11888 28364 11940 28416
rect 17224 28432 17276 28484
rect 18512 28543 18564 28552
rect 18512 28509 18521 28543
rect 18521 28509 18555 28543
rect 18555 28509 18564 28543
rect 19432 28577 19441 28611
rect 19441 28577 19475 28611
rect 19475 28577 19484 28611
rect 19432 28568 19484 28577
rect 25596 28568 25648 28620
rect 18512 28500 18564 28509
rect 18788 28500 18840 28552
rect 23388 28500 23440 28552
rect 25136 28500 25188 28552
rect 27252 28636 27304 28688
rect 29000 28636 29052 28688
rect 29552 28636 29604 28688
rect 28172 28568 28224 28620
rect 30104 28568 30156 28620
rect 31208 28611 31260 28620
rect 31208 28577 31217 28611
rect 31217 28577 31251 28611
rect 31251 28577 31260 28611
rect 31208 28568 31260 28577
rect 37188 28611 37240 28620
rect 37188 28577 37197 28611
rect 37197 28577 37231 28611
rect 37231 28577 37240 28611
rect 37188 28568 37240 28577
rect 47032 28568 47084 28620
rect 48136 28611 48188 28620
rect 48136 28577 48145 28611
rect 48145 28577 48179 28611
rect 48179 28577 48188 28611
rect 48136 28568 48188 28577
rect 20076 28432 20128 28484
rect 17684 28364 17736 28416
rect 20812 28407 20864 28416
rect 20812 28373 20821 28407
rect 20821 28373 20855 28407
rect 20855 28373 20864 28407
rect 20812 28364 20864 28373
rect 22284 28432 22336 28484
rect 23664 28432 23716 28484
rect 24032 28432 24084 28484
rect 27988 28475 28040 28484
rect 27988 28441 27997 28475
rect 27997 28441 28031 28475
rect 28031 28441 28040 28475
rect 27988 28432 28040 28441
rect 29368 28432 29420 28484
rect 30840 28500 30892 28552
rect 32772 28500 32824 28552
rect 34612 28500 34664 28552
rect 35532 28543 35584 28552
rect 35532 28509 35541 28543
rect 35541 28509 35575 28543
rect 35575 28509 35584 28543
rect 35532 28500 35584 28509
rect 34060 28432 34112 28484
rect 35716 28475 35768 28484
rect 35716 28441 35725 28475
rect 35725 28441 35759 28475
rect 35759 28441 35768 28475
rect 35716 28432 35768 28441
rect 47676 28432 47728 28484
rect 24952 28364 25004 28416
rect 25688 28407 25740 28416
rect 25688 28373 25697 28407
rect 25697 28373 25731 28407
rect 25731 28373 25740 28407
rect 25688 28364 25740 28373
rect 28356 28407 28408 28416
rect 28356 28373 28365 28407
rect 28365 28373 28399 28407
rect 28399 28373 28408 28407
rect 28356 28364 28408 28373
rect 32588 28407 32640 28416
rect 32588 28373 32597 28407
rect 32597 28373 32631 28407
rect 32631 28373 32640 28407
rect 32588 28364 32640 28373
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 8024 28160 8076 28212
rect 2872 28135 2924 28144
rect 2872 28101 2881 28135
rect 2881 28101 2915 28135
rect 2915 28101 2924 28135
rect 2872 28092 2924 28101
rect 6920 28024 6972 28076
rect 10600 28092 10652 28144
rect 12440 28160 12492 28212
rect 14280 28160 14332 28212
rect 16764 28160 16816 28212
rect 19984 28160 20036 28212
rect 23572 28160 23624 28212
rect 23664 28160 23716 28212
rect 4160 27999 4212 28008
rect 4160 27965 4169 27999
rect 4169 27965 4203 27999
rect 4203 27965 4212 27999
rect 4160 27956 4212 27965
rect 8208 28024 8260 28076
rect 9680 28024 9732 28076
rect 8944 27956 8996 28008
rect 7012 27888 7064 27940
rect 11244 27956 11296 28008
rect 11704 27956 11756 28008
rect 11796 27999 11848 28008
rect 11796 27965 11805 27999
rect 11805 27965 11839 27999
rect 11839 27965 11848 27999
rect 13820 28092 13872 28144
rect 18052 28092 18104 28144
rect 24032 28135 24084 28144
rect 24032 28101 24041 28135
rect 24041 28101 24075 28135
rect 24075 28101 24084 28135
rect 24032 28092 24084 28101
rect 25504 28160 25556 28212
rect 27712 28160 27764 28212
rect 35716 28160 35768 28212
rect 47676 28160 47728 28212
rect 47860 28160 47912 28212
rect 25136 28092 25188 28144
rect 15844 28024 15896 28076
rect 17132 28067 17184 28076
rect 17132 28033 17141 28067
rect 17141 28033 17175 28067
rect 17175 28033 17184 28067
rect 17132 28024 17184 28033
rect 18236 28067 18288 28076
rect 18236 28033 18259 28067
rect 18259 28033 18288 28067
rect 18236 28024 18288 28033
rect 14832 27999 14884 28008
rect 11796 27956 11848 27965
rect 14832 27965 14841 27999
rect 14841 27965 14875 27999
rect 14875 27965 14884 27999
rect 14832 27956 14884 27965
rect 17224 27956 17276 28008
rect 17316 27888 17368 27940
rect 18788 27956 18840 28008
rect 19156 28024 19208 28076
rect 23112 28067 23164 28076
rect 23112 28033 23121 28067
rect 23121 28033 23155 28067
rect 23155 28033 23164 28067
rect 23112 28024 23164 28033
rect 8576 27820 8628 27872
rect 24860 27956 24912 28008
rect 25688 28067 25740 28076
rect 25688 28033 25697 28067
rect 25697 28033 25731 28067
rect 25731 28033 25740 28067
rect 25688 28024 25740 28033
rect 25872 28067 25924 28076
rect 25872 28033 25881 28067
rect 25881 28033 25915 28067
rect 25915 28033 25924 28067
rect 25872 28024 25924 28033
rect 27436 28024 27488 28076
rect 26056 27956 26108 28008
rect 28356 28024 28408 28076
rect 29276 28067 29328 28076
rect 29276 28033 29285 28067
rect 29285 28033 29319 28067
rect 29319 28033 29328 28067
rect 29276 28024 29328 28033
rect 29828 28092 29880 28144
rect 34796 28092 34848 28144
rect 29644 28067 29696 28076
rect 28908 27956 28960 28008
rect 29644 28033 29653 28067
rect 29653 28033 29687 28067
rect 29687 28033 29696 28067
rect 29644 28024 29696 28033
rect 30380 28024 30432 28076
rect 32496 28024 32548 28076
rect 32772 28067 32824 28076
rect 32772 28033 32781 28067
rect 32781 28033 32815 28067
rect 32815 28033 32824 28067
rect 32772 28024 32824 28033
rect 33416 28024 33468 28076
rect 37280 28067 37332 28076
rect 37280 28033 37289 28067
rect 37289 28033 37323 28067
rect 37323 28033 37332 28067
rect 37280 28024 37332 28033
rect 47860 28067 47912 28076
rect 47860 28033 47869 28067
rect 47869 28033 47903 28067
rect 47903 28033 47912 28067
rect 47860 28024 47912 28033
rect 30748 27956 30800 28008
rect 31300 27956 31352 28008
rect 33232 27999 33284 28008
rect 33232 27965 33241 27999
rect 33241 27965 33275 27999
rect 33275 27965 33284 27999
rect 33232 27956 33284 27965
rect 36452 27956 36504 28008
rect 27896 27888 27948 27940
rect 35532 27888 35584 27940
rect 19432 27820 19484 27872
rect 19708 27820 19760 27872
rect 20444 27863 20496 27872
rect 20444 27829 20453 27863
rect 20453 27829 20487 27863
rect 20487 27829 20496 27863
rect 20444 27820 20496 27829
rect 22744 27820 22796 27872
rect 25320 27820 25372 27872
rect 27344 27863 27396 27872
rect 27344 27829 27353 27863
rect 27353 27829 27387 27863
rect 27387 27829 27396 27863
rect 27344 27820 27396 27829
rect 29000 27863 29052 27872
rect 29000 27829 29009 27863
rect 29009 27829 29043 27863
rect 29043 27829 29052 27863
rect 29000 27820 29052 27829
rect 48044 27863 48096 27872
rect 48044 27829 48053 27863
rect 48053 27829 48087 27863
rect 48087 27829 48096 27863
rect 48044 27820 48096 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 17224 27659 17276 27668
rect 8944 27591 8996 27600
rect 8944 27557 8953 27591
rect 8953 27557 8987 27591
rect 8987 27557 8996 27591
rect 8944 27548 8996 27557
rect 17224 27625 17233 27659
rect 17233 27625 17267 27659
rect 17267 27625 17276 27659
rect 17224 27616 17276 27625
rect 11152 27591 11204 27600
rect 1400 27412 1452 27464
rect 2228 27412 2280 27464
rect 1768 27344 1820 27396
rect 6920 27412 6972 27464
rect 8484 27412 8536 27464
rect 3332 27344 3384 27396
rect 11152 27557 11161 27591
rect 11161 27557 11195 27591
rect 11195 27557 11204 27591
rect 11152 27548 11204 27557
rect 11244 27548 11296 27600
rect 13084 27548 13136 27600
rect 16120 27548 16172 27600
rect 16672 27548 16724 27600
rect 9128 27480 9180 27532
rect 9680 27480 9732 27532
rect 15752 27480 15804 27532
rect 16580 27523 16632 27532
rect 16580 27489 16589 27523
rect 16589 27489 16623 27523
rect 16623 27489 16632 27523
rect 16580 27480 16632 27489
rect 20076 27616 20128 27668
rect 24952 27616 25004 27668
rect 25688 27616 25740 27668
rect 21088 27591 21140 27600
rect 21088 27557 21097 27591
rect 21097 27557 21131 27591
rect 21131 27557 21140 27591
rect 21088 27548 21140 27557
rect 22560 27548 22612 27600
rect 34612 27616 34664 27668
rect 34336 27548 34388 27600
rect 47308 27548 47360 27600
rect 9588 27455 9640 27464
rect 1952 27276 2004 27328
rect 8208 27319 8260 27328
rect 8208 27285 8217 27319
rect 8217 27285 8251 27319
rect 8251 27285 8260 27319
rect 8208 27276 8260 27285
rect 9588 27421 9597 27455
rect 9597 27421 9631 27455
rect 9631 27421 9640 27455
rect 9588 27412 9640 27421
rect 11888 27455 11940 27464
rect 9496 27344 9548 27396
rect 10784 27387 10836 27396
rect 10784 27353 10793 27387
rect 10793 27353 10827 27387
rect 10827 27353 10836 27387
rect 10784 27344 10836 27353
rect 11888 27421 11922 27455
rect 11922 27421 11940 27455
rect 11888 27412 11940 27421
rect 16396 27412 16448 27464
rect 17132 27455 17184 27464
rect 11796 27344 11848 27396
rect 17132 27421 17141 27455
rect 17141 27421 17175 27455
rect 17175 27421 17184 27455
rect 17132 27412 17184 27421
rect 17316 27412 17368 27464
rect 9772 27276 9824 27328
rect 10232 27276 10284 27328
rect 11060 27276 11112 27328
rect 11244 27276 11296 27328
rect 13268 27276 13320 27328
rect 14280 27276 14332 27328
rect 16304 27276 16356 27328
rect 18696 27455 18748 27464
rect 18696 27421 18705 27455
rect 18705 27421 18739 27455
rect 18739 27421 18748 27455
rect 18696 27412 18748 27421
rect 19708 27455 19760 27464
rect 19708 27421 19717 27455
rect 19717 27421 19751 27455
rect 19751 27421 19760 27455
rect 19708 27412 19760 27421
rect 25780 27480 25832 27532
rect 26792 27523 26844 27532
rect 26792 27489 26801 27523
rect 26801 27489 26835 27523
rect 26835 27489 26844 27523
rect 26792 27480 26844 27489
rect 29552 27523 29604 27532
rect 29552 27489 29561 27523
rect 29561 27489 29595 27523
rect 29595 27489 29604 27523
rect 29552 27480 29604 27489
rect 30564 27480 30616 27532
rect 37096 27523 37148 27532
rect 37096 27489 37105 27523
rect 37105 27489 37139 27523
rect 37139 27489 37148 27523
rect 37096 27480 37148 27489
rect 19340 27344 19392 27396
rect 19984 27387 20036 27396
rect 19984 27353 20018 27387
rect 20018 27353 20036 27387
rect 19984 27344 20036 27353
rect 21272 27344 21324 27396
rect 23664 27412 23716 27464
rect 24952 27455 25004 27464
rect 24952 27421 24961 27455
rect 24961 27421 24995 27455
rect 24995 27421 25004 27455
rect 24952 27412 25004 27421
rect 27252 27455 27304 27464
rect 27252 27421 27261 27455
rect 27261 27421 27295 27455
rect 27295 27421 27304 27455
rect 27252 27412 27304 27421
rect 27344 27412 27396 27464
rect 29000 27412 29052 27464
rect 32772 27412 32824 27464
rect 34704 27455 34756 27464
rect 34704 27421 34713 27455
rect 34713 27421 34747 27455
rect 34747 27421 34756 27455
rect 34704 27412 34756 27421
rect 47308 27412 47360 27464
rect 47676 27412 47728 27464
rect 22468 27276 22520 27328
rect 22560 27276 22612 27328
rect 23020 27276 23072 27328
rect 28632 27319 28684 27328
rect 28632 27285 28641 27319
rect 28641 27285 28675 27319
rect 28675 27285 28684 27319
rect 28632 27276 28684 27285
rect 29184 27276 29236 27328
rect 33508 27344 33560 27396
rect 37372 27344 37424 27396
rect 33600 27276 33652 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 9404 27072 9456 27124
rect 9588 27072 9640 27124
rect 13084 27072 13136 27124
rect 13268 27072 13320 27124
rect 14372 27072 14424 27124
rect 14832 27072 14884 27124
rect 15016 27072 15068 27124
rect 15660 27072 15712 27124
rect 1952 27047 2004 27056
rect 1952 27013 1961 27047
rect 1961 27013 1995 27047
rect 1995 27013 2004 27047
rect 1952 27004 2004 27013
rect 6552 27004 6604 27056
rect 1768 26979 1820 26988
rect 1768 26945 1777 26979
rect 1777 26945 1811 26979
rect 1811 26945 1820 26979
rect 1768 26936 1820 26945
rect 7196 26936 7248 26988
rect 8024 26936 8076 26988
rect 2780 26911 2832 26920
rect 2780 26877 2789 26911
rect 2789 26877 2823 26911
rect 2823 26877 2832 26911
rect 2780 26868 2832 26877
rect 7380 26868 7432 26920
rect 8208 26868 8260 26920
rect 10784 26936 10836 26988
rect 12624 26936 12676 26988
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 13820 26936 13872 26945
rect 15016 26936 15068 26988
rect 15752 26979 15804 26988
rect 15752 26945 15761 26979
rect 15761 26945 15795 26979
rect 15795 26945 15804 26979
rect 15752 26936 15804 26945
rect 16672 26936 16724 26988
rect 14096 26868 14148 26920
rect 14188 26868 14240 26920
rect 16396 26868 16448 26920
rect 17500 27004 17552 27056
rect 17040 26936 17092 26988
rect 17408 26979 17460 26988
rect 17408 26945 17417 26979
rect 17417 26945 17451 26979
rect 17451 26945 17460 26979
rect 18512 27072 18564 27124
rect 19340 27072 19392 27124
rect 20260 27072 20312 27124
rect 24952 27072 25004 27124
rect 25044 27072 25096 27124
rect 17868 27004 17920 27056
rect 17408 26936 17460 26945
rect 18788 26936 18840 26988
rect 20812 27004 20864 27056
rect 22744 27047 22796 27056
rect 22744 27013 22753 27047
rect 22753 27013 22787 27047
rect 22787 27013 22796 27047
rect 22744 27004 22796 27013
rect 25320 27047 25372 27056
rect 25320 27013 25354 27047
rect 25354 27013 25372 27047
rect 25320 27004 25372 27013
rect 28908 27004 28960 27056
rect 29184 27047 29236 27056
rect 29184 27013 29193 27047
rect 29193 27013 29227 27047
rect 29227 27013 29236 27047
rect 29184 27004 29236 27013
rect 29644 27072 29696 27124
rect 32128 27072 32180 27124
rect 34704 27072 34756 27124
rect 37372 27115 37424 27124
rect 30564 27004 30616 27056
rect 32588 27004 32640 27056
rect 33692 27004 33744 27056
rect 20444 26936 20496 26988
rect 22560 26979 22612 26988
rect 22560 26945 22569 26979
rect 22569 26945 22603 26979
rect 22603 26945 22612 26979
rect 22560 26936 22612 26945
rect 26332 26936 26384 26988
rect 27252 26936 27304 26988
rect 27436 26979 27488 26988
rect 27436 26945 27445 26979
rect 27445 26945 27479 26979
rect 27479 26945 27488 26979
rect 27436 26936 27488 26945
rect 28172 26936 28224 26988
rect 29368 26979 29420 26988
rect 29368 26945 29377 26979
rect 29377 26945 29411 26979
rect 29411 26945 29420 26979
rect 29368 26936 29420 26945
rect 30380 26936 30432 26988
rect 32220 26936 32272 26988
rect 14280 26800 14332 26852
rect 15752 26800 15804 26852
rect 16304 26800 16356 26852
rect 18512 26800 18564 26852
rect 6736 26732 6788 26784
rect 13820 26732 13872 26784
rect 16764 26732 16816 26784
rect 23756 26868 23808 26920
rect 23940 26911 23992 26920
rect 23940 26877 23949 26911
rect 23949 26877 23983 26911
rect 23983 26877 23992 26911
rect 23940 26868 23992 26877
rect 26424 26868 26476 26920
rect 18880 26800 18932 26852
rect 19432 26800 19484 26852
rect 20444 26732 20496 26784
rect 24952 26732 25004 26784
rect 29552 26800 29604 26852
rect 30472 26868 30524 26920
rect 31484 26868 31536 26920
rect 32496 26868 32548 26920
rect 34796 26936 34848 26988
rect 35808 26936 35860 26988
rect 37372 27081 37381 27115
rect 37381 27081 37415 27115
rect 37415 27081 37424 27115
rect 37372 27072 37424 27081
rect 37280 26979 37332 26988
rect 37280 26945 37289 26979
rect 37289 26945 37323 26979
rect 37323 26945 37332 26979
rect 37280 26936 37332 26945
rect 34704 26911 34756 26920
rect 34704 26877 34713 26911
rect 34713 26877 34747 26911
rect 34747 26877 34756 26911
rect 34704 26868 34756 26877
rect 33324 26800 33376 26852
rect 26056 26732 26108 26784
rect 26700 26732 26752 26784
rect 26884 26732 26936 26784
rect 27252 26732 27304 26784
rect 27620 26732 27672 26784
rect 29644 26732 29696 26784
rect 36268 26732 36320 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 3792 26528 3844 26580
rect 15660 26528 15712 26580
rect 15752 26528 15804 26580
rect 4804 26460 4856 26512
rect 14740 26503 14792 26512
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 2780 26435 2832 26444
rect 2780 26401 2789 26435
rect 2789 26401 2823 26435
rect 2823 26401 2832 26435
rect 6552 26435 6604 26444
rect 2780 26392 2832 26401
rect 6552 26401 6561 26435
rect 6561 26401 6595 26435
rect 6595 26401 6604 26435
rect 6552 26392 6604 26401
rect 6736 26435 6788 26444
rect 6736 26401 6745 26435
rect 6745 26401 6779 26435
rect 6779 26401 6788 26435
rect 6736 26392 6788 26401
rect 1584 26299 1636 26308
rect 1584 26265 1593 26299
rect 1593 26265 1627 26299
rect 1627 26265 1636 26299
rect 1584 26256 1636 26265
rect 3976 26256 4028 26308
rect 8576 26392 8628 26444
rect 10508 26435 10560 26444
rect 10508 26401 10517 26435
rect 10517 26401 10551 26435
rect 10551 26401 10560 26435
rect 10508 26392 10560 26401
rect 14740 26469 14749 26503
rect 14749 26469 14783 26503
rect 14783 26469 14792 26503
rect 14740 26460 14792 26469
rect 16672 26528 16724 26580
rect 17040 26528 17092 26580
rect 17408 26528 17460 26580
rect 18512 26528 18564 26580
rect 30840 26528 30892 26580
rect 46572 26528 46624 26580
rect 17500 26460 17552 26512
rect 17684 26460 17736 26512
rect 24032 26460 24084 26512
rect 25228 26460 25280 26512
rect 25872 26460 25924 26512
rect 9128 26299 9180 26308
rect 9128 26265 9137 26299
rect 9137 26265 9171 26299
rect 9171 26265 9180 26299
rect 9128 26256 9180 26265
rect 13268 26256 13320 26308
rect 15384 26367 15436 26376
rect 15384 26333 15393 26367
rect 15393 26333 15427 26367
rect 15427 26333 15436 26367
rect 15384 26324 15436 26333
rect 16396 26324 16448 26376
rect 15476 26256 15528 26308
rect 16672 26256 16724 26308
rect 17132 26324 17184 26376
rect 18604 26324 18656 26376
rect 19432 26324 19484 26376
rect 20628 26324 20680 26376
rect 23020 26324 23072 26376
rect 26056 26392 26108 26444
rect 26240 26392 26292 26444
rect 26148 26367 26200 26376
rect 26148 26333 26157 26367
rect 26157 26333 26191 26367
rect 26191 26333 26200 26367
rect 26148 26324 26200 26333
rect 27252 26367 27304 26376
rect 23664 26299 23716 26308
rect 23664 26265 23673 26299
rect 23673 26265 23707 26299
rect 23707 26265 23716 26299
rect 23664 26256 23716 26265
rect 24768 26256 24820 26308
rect 24952 26256 25004 26308
rect 25688 26256 25740 26308
rect 27252 26333 27261 26367
rect 27261 26333 27295 26367
rect 27295 26333 27304 26367
rect 27252 26324 27304 26333
rect 45744 26460 45796 26512
rect 30840 26435 30892 26444
rect 30840 26401 30849 26435
rect 30849 26401 30883 26435
rect 30883 26401 30892 26435
rect 30840 26392 30892 26401
rect 32404 26435 32456 26444
rect 32404 26401 32413 26435
rect 32413 26401 32447 26435
rect 32447 26401 32456 26435
rect 32404 26392 32456 26401
rect 33600 26392 33652 26444
rect 36268 26392 36320 26444
rect 28448 26367 28500 26376
rect 28448 26333 28457 26367
rect 28457 26333 28491 26367
rect 28491 26333 28500 26367
rect 28448 26324 28500 26333
rect 31944 26324 31996 26376
rect 26424 26256 26476 26308
rect 2228 26188 2280 26240
rect 17316 26188 17368 26240
rect 18236 26188 18288 26240
rect 19248 26188 19300 26240
rect 20444 26188 20496 26240
rect 23388 26188 23440 26240
rect 24032 26188 24084 26240
rect 27344 26231 27396 26240
rect 27344 26197 27353 26231
rect 27353 26197 27387 26231
rect 27387 26197 27396 26231
rect 27344 26188 27396 26197
rect 30380 26256 30432 26308
rect 30472 26188 30524 26240
rect 34796 26324 34848 26376
rect 33968 26256 34020 26308
rect 45928 26392 45980 26444
rect 44824 26256 44876 26308
rect 47952 26299 48004 26308
rect 47952 26265 47961 26299
rect 47961 26265 47995 26299
rect 47995 26265 48004 26299
rect 47952 26256 48004 26265
rect 48136 26299 48188 26308
rect 48136 26265 48145 26299
rect 48145 26265 48179 26299
rect 48179 26265 48188 26299
rect 48136 26256 48188 26265
rect 35164 26188 35216 26240
rect 35808 26188 35860 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 1584 25984 1636 26036
rect 2964 25984 3016 26036
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 2228 25891 2280 25900
rect 2228 25857 2237 25891
rect 2237 25857 2271 25891
rect 2271 25857 2280 25891
rect 2228 25848 2280 25857
rect 6644 25891 6696 25900
rect 6644 25857 6653 25891
rect 6653 25857 6687 25891
rect 6687 25857 6696 25891
rect 6644 25848 6696 25857
rect 6276 25780 6328 25832
rect 6828 25687 6880 25696
rect 6828 25653 6837 25687
rect 6837 25653 6871 25687
rect 6871 25653 6880 25687
rect 6828 25644 6880 25653
rect 9128 25984 9180 26036
rect 16672 26027 16724 26036
rect 16672 25993 16681 26027
rect 16681 25993 16715 26027
rect 16715 25993 16724 26027
rect 16672 25984 16724 25993
rect 17040 26027 17092 26036
rect 17040 25993 17049 26027
rect 17049 25993 17083 26027
rect 17083 25993 17092 26027
rect 17040 25984 17092 25993
rect 25228 25984 25280 26036
rect 7748 25848 7800 25900
rect 17408 25916 17460 25968
rect 26056 25916 26108 25968
rect 28172 25984 28224 26036
rect 28448 25984 28500 26036
rect 26976 25916 27028 25968
rect 28356 25916 28408 25968
rect 8300 25848 8352 25900
rect 9312 25891 9364 25900
rect 9312 25857 9321 25891
rect 9321 25857 9355 25891
rect 9355 25857 9364 25891
rect 9312 25848 9364 25857
rect 10232 25848 10284 25900
rect 13268 25891 13320 25900
rect 9220 25780 9272 25832
rect 11612 25823 11664 25832
rect 11612 25789 11621 25823
rect 11621 25789 11655 25823
rect 11655 25789 11664 25823
rect 11612 25780 11664 25789
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 14188 25891 14240 25900
rect 14188 25857 14197 25891
rect 14197 25857 14231 25891
rect 14231 25857 14240 25891
rect 14188 25848 14240 25857
rect 16948 25848 17000 25900
rect 17132 25891 17184 25900
rect 17132 25857 17141 25891
rect 17141 25857 17175 25891
rect 17175 25857 17184 25891
rect 17132 25848 17184 25857
rect 14280 25823 14332 25832
rect 14280 25789 14289 25823
rect 14289 25789 14323 25823
rect 14323 25789 14332 25823
rect 14280 25780 14332 25789
rect 18236 25823 18288 25832
rect 18236 25789 18245 25823
rect 18245 25789 18279 25823
rect 18279 25789 18288 25823
rect 18236 25780 18288 25789
rect 19524 25780 19576 25832
rect 12716 25712 12768 25764
rect 19248 25712 19300 25764
rect 23480 25891 23532 25900
rect 23480 25857 23489 25891
rect 23489 25857 23523 25891
rect 23523 25857 23532 25891
rect 23480 25848 23532 25857
rect 24584 25891 24636 25900
rect 23572 25823 23624 25832
rect 23572 25789 23581 25823
rect 23581 25789 23615 25823
rect 23615 25789 23624 25823
rect 23572 25780 23624 25789
rect 24584 25857 24593 25891
rect 24593 25857 24627 25891
rect 24627 25857 24636 25891
rect 24584 25848 24636 25857
rect 26148 25848 26200 25900
rect 29644 25959 29696 25968
rect 29644 25925 29653 25959
rect 29653 25925 29687 25959
rect 29687 25925 29696 25959
rect 29644 25916 29696 25925
rect 29184 25848 29236 25900
rect 32036 25916 32088 25968
rect 32496 25848 32548 25900
rect 20444 25712 20496 25764
rect 22376 25712 22428 25764
rect 24860 25712 24912 25764
rect 10968 25644 11020 25696
rect 12072 25644 12124 25696
rect 12256 25644 12308 25696
rect 16948 25644 17000 25696
rect 17408 25644 17460 25696
rect 18236 25644 18288 25696
rect 19432 25644 19484 25696
rect 19616 25687 19668 25696
rect 19616 25653 19625 25687
rect 19625 25653 19659 25687
rect 19659 25653 19668 25687
rect 19616 25644 19668 25653
rect 19708 25644 19760 25696
rect 23940 25687 23992 25696
rect 23940 25653 23949 25687
rect 23949 25653 23983 25687
rect 23983 25653 23992 25687
rect 23940 25644 23992 25653
rect 25136 25823 25188 25832
rect 25136 25789 25145 25823
rect 25145 25789 25179 25823
rect 25179 25789 25188 25823
rect 25136 25780 25188 25789
rect 25504 25780 25556 25832
rect 31024 25823 31076 25832
rect 31024 25789 31033 25823
rect 31033 25789 31067 25823
rect 31067 25789 31076 25823
rect 31024 25780 31076 25789
rect 31576 25780 31628 25832
rect 33048 25823 33100 25832
rect 33048 25789 33057 25823
rect 33057 25789 33091 25823
rect 33091 25789 33100 25823
rect 33048 25780 33100 25789
rect 45560 25916 45612 25968
rect 35164 25891 35216 25900
rect 35164 25857 35173 25891
rect 35173 25857 35207 25891
rect 35207 25857 35216 25891
rect 35164 25848 35216 25857
rect 35808 25823 35860 25832
rect 35808 25789 35817 25823
rect 35817 25789 35851 25823
rect 35851 25789 35860 25823
rect 35808 25780 35860 25789
rect 46664 25780 46716 25832
rect 25228 25712 25280 25764
rect 33968 25712 34020 25764
rect 27160 25644 27212 25696
rect 27988 25644 28040 25696
rect 31944 25644 31996 25696
rect 32496 25644 32548 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6828 25440 6880 25492
rect 19708 25440 19760 25492
rect 23204 25483 23256 25492
rect 9220 25347 9272 25356
rect 9220 25313 9229 25347
rect 9229 25313 9263 25347
rect 9263 25313 9272 25347
rect 9220 25304 9272 25313
rect 9772 25372 9824 25424
rect 10784 25372 10836 25424
rect 11336 25372 11388 25424
rect 12072 25415 12124 25424
rect 12072 25381 12081 25415
rect 12081 25381 12115 25415
rect 12115 25381 12124 25415
rect 12072 25372 12124 25381
rect 13176 25372 13228 25424
rect 9864 25304 9916 25356
rect 8760 25236 8812 25288
rect 9588 25279 9640 25288
rect 9588 25245 9597 25279
rect 9597 25245 9631 25279
rect 9631 25245 9640 25279
rect 9588 25236 9640 25245
rect 8300 25168 8352 25220
rect 10784 25279 10836 25288
rect 10784 25245 10793 25279
rect 10793 25245 10827 25279
rect 10827 25245 10836 25279
rect 10784 25236 10836 25245
rect 10876 25279 10928 25288
rect 10876 25245 10885 25279
rect 10885 25245 10919 25279
rect 10919 25245 10928 25279
rect 12992 25304 13044 25356
rect 14464 25372 14516 25424
rect 17316 25372 17368 25424
rect 23204 25449 23213 25483
rect 23213 25449 23247 25483
rect 23247 25449 23256 25483
rect 23204 25440 23256 25449
rect 23572 25483 23624 25492
rect 23572 25449 23581 25483
rect 23581 25449 23615 25483
rect 23615 25449 23624 25483
rect 23572 25440 23624 25449
rect 25136 25440 25188 25492
rect 26148 25440 26200 25492
rect 24492 25372 24544 25424
rect 24860 25372 24912 25424
rect 28356 25440 28408 25492
rect 28816 25440 28868 25492
rect 30932 25440 30984 25492
rect 47124 25440 47176 25492
rect 27160 25372 27212 25424
rect 38476 25372 38528 25424
rect 13452 25304 13504 25356
rect 10876 25236 10928 25245
rect 12256 25279 12308 25288
rect 12256 25245 12265 25279
rect 12265 25245 12299 25279
rect 12299 25245 12308 25279
rect 12256 25236 12308 25245
rect 13912 25236 13964 25288
rect 14188 25236 14240 25288
rect 14464 25279 14516 25288
rect 14464 25245 14473 25279
rect 14473 25245 14507 25279
rect 14507 25245 14516 25279
rect 14464 25236 14516 25245
rect 15384 25304 15436 25356
rect 16212 25347 16264 25356
rect 16212 25313 16221 25347
rect 16221 25313 16255 25347
rect 16255 25313 16264 25347
rect 16212 25304 16264 25313
rect 16764 25236 16816 25288
rect 17040 25236 17092 25288
rect 19156 25236 19208 25288
rect 19432 25304 19484 25356
rect 20076 25304 20128 25356
rect 21548 25304 21600 25356
rect 19524 25279 19576 25288
rect 19524 25245 19533 25279
rect 19533 25245 19567 25279
rect 19567 25245 19576 25279
rect 19524 25236 19576 25245
rect 24584 25279 24636 25288
rect 2044 25100 2096 25152
rect 9128 25100 9180 25152
rect 9312 25100 9364 25152
rect 20812 25211 20864 25220
rect 20812 25177 20846 25211
rect 20846 25177 20864 25211
rect 20812 25168 20864 25177
rect 13544 25143 13596 25152
rect 13544 25109 13553 25143
rect 13553 25109 13587 25143
rect 13587 25109 13596 25143
rect 13544 25100 13596 25109
rect 14372 25143 14424 25152
rect 14372 25109 14381 25143
rect 14381 25109 14415 25143
rect 14415 25109 14424 25143
rect 14372 25100 14424 25109
rect 16580 25100 16632 25152
rect 19156 25100 19208 25152
rect 19340 25100 19392 25152
rect 19984 25100 20036 25152
rect 21548 25100 21600 25152
rect 22192 25168 22244 25220
rect 23204 25168 23256 25220
rect 24584 25245 24593 25279
rect 24593 25245 24627 25279
rect 24627 25245 24636 25279
rect 24584 25236 24636 25245
rect 26148 25279 26200 25288
rect 26148 25245 26157 25279
rect 26157 25245 26191 25279
rect 26191 25245 26200 25279
rect 26148 25236 26200 25245
rect 27988 25279 28040 25288
rect 27988 25245 27997 25279
rect 27997 25245 28031 25279
rect 28031 25245 28040 25279
rect 27988 25236 28040 25245
rect 29644 25236 29696 25288
rect 26240 25168 26292 25220
rect 27436 25168 27488 25220
rect 28264 25168 28316 25220
rect 28816 25211 28868 25220
rect 28816 25177 28825 25211
rect 28825 25177 28859 25211
rect 28859 25177 28868 25211
rect 28816 25168 28868 25177
rect 28908 25168 28960 25220
rect 33508 25304 33560 25356
rect 32496 25236 32548 25288
rect 33692 25236 33744 25288
rect 47860 25279 47912 25288
rect 47860 25245 47869 25279
rect 47869 25245 47903 25279
rect 47903 25245 47912 25279
rect 47860 25236 47912 25245
rect 26976 25100 27028 25152
rect 30932 25100 30984 25152
rect 40132 25168 40184 25220
rect 33508 25100 33560 25152
rect 33692 25100 33744 25152
rect 34796 25143 34848 25152
rect 34796 25109 34805 25143
rect 34805 25109 34839 25143
rect 34839 25109 34848 25143
rect 34796 25100 34848 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 9404 24828 9456 24880
rect 7564 24803 7616 24812
rect 7564 24769 7573 24803
rect 7573 24769 7607 24803
rect 7607 24769 7616 24803
rect 7564 24760 7616 24769
rect 7656 24760 7708 24812
rect 8392 24803 8444 24812
rect 8392 24769 8401 24803
rect 8401 24769 8435 24803
rect 8435 24769 8444 24803
rect 8392 24760 8444 24769
rect 8760 24735 8812 24744
rect 8760 24701 8769 24735
rect 8769 24701 8803 24735
rect 8803 24701 8812 24735
rect 8760 24692 8812 24701
rect 9220 24760 9272 24812
rect 9677 24803 9729 24812
rect 9677 24769 9704 24803
rect 9704 24769 9729 24803
rect 9677 24760 9729 24769
rect 9956 24803 10008 24812
rect 9956 24769 9965 24803
rect 9965 24769 9999 24803
rect 9999 24769 10008 24803
rect 11980 24896 12032 24948
rect 23480 24939 23532 24948
rect 10968 24828 11020 24880
rect 19984 24828 20036 24880
rect 23480 24905 23489 24939
rect 23489 24905 23523 24939
rect 23523 24905 23532 24939
rect 23480 24896 23532 24905
rect 24032 24828 24084 24880
rect 26976 24896 27028 24948
rect 48044 24896 48096 24948
rect 9956 24760 10008 24769
rect 10324 24692 10376 24744
rect 11612 24692 11664 24744
rect 13176 24760 13228 24812
rect 16580 24760 16632 24812
rect 18880 24760 18932 24812
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 19340 24803 19392 24812
rect 19340 24769 19349 24803
rect 19349 24769 19383 24803
rect 19383 24769 19392 24803
rect 19340 24760 19392 24769
rect 19892 24760 19944 24812
rect 20803 24809 20855 24812
rect 20803 24775 20836 24809
rect 20836 24775 20855 24809
rect 20803 24760 20855 24775
rect 21180 24760 21232 24812
rect 21364 24760 21416 24812
rect 14372 24692 14424 24744
rect 20076 24692 20128 24744
rect 20996 24692 21048 24744
rect 2228 24556 2280 24608
rect 8668 24599 8720 24608
rect 8668 24565 8677 24599
rect 8677 24565 8711 24599
rect 8711 24565 8720 24599
rect 8668 24556 8720 24565
rect 9220 24556 9272 24608
rect 10876 24556 10928 24608
rect 13452 24556 13504 24608
rect 14280 24556 14332 24608
rect 15108 24556 15160 24608
rect 20352 24624 20404 24676
rect 20628 24624 20680 24676
rect 21640 24624 21692 24676
rect 18880 24556 18932 24608
rect 22928 24556 22980 24608
rect 23756 24760 23808 24812
rect 32036 24828 32088 24880
rect 33048 24828 33100 24880
rect 25688 24803 25740 24812
rect 24124 24692 24176 24744
rect 25688 24769 25697 24803
rect 25697 24769 25731 24803
rect 25731 24769 25740 24803
rect 25688 24760 25740 24769
rect 25872 24803 25924 24812
rect 25872 24769 25881 24803
rect 25881 24769 25915 24803
rect 25915 24769 25924 24803
rect 25872 24760 25924 24769
rect 27344 24760 27396 24812
rect 27988 24760 28040 24812
rect 31944 24760 31996 24812
rect 32496 24760 32548 24812
rect 38016 24803 38068 24812
rect 38016 24769 38025 24803
rect 38025 24769 38059 24803
rect 38059 24769 38068 24803
rect 38016 24760 38068 24769
rect 38292 24803 38344 24812
rect 38292 24769 38301 24803
rect 38301 24769 38335 24803
rect 38335 24769 38344 24803
rect 38292 24760 38344 24769
rect 45652 24760 45704 24812
rect 47216 24760 47268 24812
rect 27160 24692 27212 24744
rect 29552 24692 29604 24744
rect 31392 24692 31444 24744
rect 32588 24692 32640 24744
rect 32956 24735 33008 24744
rect 32956 24701 32965 24735
rect 32965 24701 32999 24735
rect 32999 24701 33008 24735
rect 32956 24692 33008 24701
rect 34428 24735 34480 24744
rect 34428 24701 34437 24735
rect 34437 24701 34471 24735
rect 34471 24701 34480 24735
rect 34428 24692 34480 24701
rect 38108 24735 38160 24744
rect 38108 24701 38117 24735
rect 38117 24701 38151 24735
rect 38151 24701 38160 24735
rect 38108 24692 38160 24701
rect 40040 24735 40092 24744
rect 40040 24701 40049 24735
rect 40049 24701 40083 24735
rect 40083 24701 40092 24735
rect 40040 24692 40092 24701
rect 40224 24735 40276 24744
rect 40224 24701 40233 24735
rect 40233 24701 40267 24735
rect 40267 24701 40276 24735
rect 40224 24692 40276 24701
rect 41236 24735 41288 24744
rect 41236 24701 41245 24735
rect 41245 24701 41279 24735
rect 41279 24701 41288 24735
rect 41236 24692 41288 24701
rect 23204 24556 23256 24608
rect 23388 24556 23440 24608
rect 23664 24556 23716 24608
rect 24768 24556 24820 24608
rect 25872 24556 25924 24608
rect 26424 24556 26476 24608
rect 27988 24556 28040 24608
rect 29736 24556 29788 24608
rect 35624 24556 35676 24608
rect 38108 24599 38160 24608
rect 38108 24565 38117 24599
rect 38117 24565 38151 24599
rect 38151 24565 38160 24599
rect 38108 24556 38160 24565
rect 38476 24599 38528 24608
rect 38476 24565 38485 24599
rect 38485 24565 38519 24599
rect 38519 24565 38528 24599
rect 38476 24556 38528 24565
rect 38660 24624 38712 24676
rect 48136 24624 48188 24676
rect 44916 24556 44968 24608
rect 46296 24556 46348 24608
rect 47676 24599 47728 24608
rect 47676 24565 47685 24599
rect 47685 24565 47719 24599
rect 47719 24565 47728 24599
rect 47676 24556 47728 24565
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 8392 24352 8444 24404
rect 9956 24352 10008 24404
rect 10416 24352 10468 24404
rect 12900 24395 12952 24404
rect 12900 24361 12909 24395
rect 12909 24361 12943 24395
rect 12943 24361 12952 24395
rect 12900 24352 12952 24361
rect 7564 24284 7616 24336
rect 9588 24216 9640 24268
rect 10324 24216 10376 24268
rect 19432 24216 19484 24268
rect 1400 24191 1452 24200
rect 1400 24157 1409 24191
rect 1409 24157 1443 24191
rect 1443 24157 1452 24191
rect 1400 24148 1452 24157
rect 9036 24191 9088 24200
rect 9036 24157 9045 24191
rect 9045 24157 9079 24191
rect 9079 24157 9088 24191
rect 9036 24148 9088 24157
rect 9680 24191 9732 24200
rect 7656 24080 7708 24132
rect 9680 24157 9689 24191
rect 9689 24157 9723 24191
rect 9723 24157 9732 24191
rect 9680 24148 9732 24157
rect 22744 24352 22796 24404
rect 22836 24352 22888 24404
rect 24308 24352 24360 24404
rect 23020 24284 23072 24336
rect 38660 24352 38712 24404
rect 40224 24395 40276 24404
rect 40224 24361 40233 24395
rect 40233 24361 40267 24395
rect 40267 24361 40276 24395
rect 40224 24352 40276 24361
rect 32496 24284 32548 24336
rect 33692 24284 33744 24336
rect 34796 24284 34848 24336
rect 23940 24216 23992 24268
rect 24492 24259 24544 24268
rect 24492 24225 24501 24259
rect 24501 24225 24535 24259
rect 24535 24225 24544 24259
rect 24492 24216 24544 24225
rect 29092 24216 29144 24268
rect 35624 24284 35676 24336
rect 48044 24284 48096 24336
rect 36544 24259 36596 24268
rect 36544 24225 36553 24259
rect 36553 24225 36587 24259
rect 36587 24225 36596 24259
rect 36544 24216 36596 24225
rect 46296 24259 46348 24268
rect 46296 24225 46305 24259
rect 46305 24225 46339 24259
rect 46339 24225 46348 24259
rect 46296 24216 46348 24225
rect 47676 24216 47728 24268
rect 48136 24259 48188 24268
rect 48136 24225 48145 24259
rect 48145 24225 48179 24259
rect 48179 24225 48188 24259
rect 48136 24216 48188 24225
rect 10048 24080 10100 24132
rect 1584 24055 1636 24064
rect 1584 24021 1593 24055
rect 1593 24021 1627 24055
rect 1627 24021 1636 24055
rect 1584 24012 1636 24021
rect 7288 24012 7340 24064
rect 21824 24148 21876 24200
rect 24400 24191 24452 24200
rect 24400 24157 24409 24191
rect 24409 24157 24443 24191
rect 24443 24157 24452 24191
rect 24676 24191 24728 24200
rect 24400 24148 24452 24157
rect 24676 24157 24685 24191
rect 24685 24157 24719 24191
rect 24719 24157 24728 24191
rect 24676 24148 24728 24157
rect 27620 24191 27672 24200
rect 27620 24157 27629 24191
rect 27629 24157 27663 24191
rect 27663 24157 27672 24191
rect 27620 24148 27672 24157
rect 12532 24080 12584 24132
rect 13268 24080 13320 24132
rect 16580 24123 16632 24132
rect 12808 24012 12860 24064
rect 13084 24055 13136 24064
rect 13084 24021 13093 24055
rect 13093 24021 13127 24055
rect 13127 24021 13136 24055
rect 13084 24012 13136 24021
rect 16580 24089 16589 24123
rect 16589 24089 16623 24123
rect 16623 24089 16632 24123
rect 16580 24080 16632 24089
rect 17960 24080 18012 24132
rect 20352 24080 20404 24132
rect 21640 24123 21692 24132
rect 21640 24089 21649 24123
rect 21649 24089 21683 24123
rect 21683 24089 21692 24123
rect 21640 24080 21692 24089
rect 21732 24080 21784 24132
rect 17132 24012 17184 24064
rect 17224 24012 17276 24064
rect 20628 24012 20680 24064
rect 20720 24012 20772 24064
rect 22744 24080 22796 24132
rect 25872 24080 25924 24132
rect 27896 24123 27948 24132
rect 27896 24089 27930 24123
rect 27930 24089 27948 24123
rect 28172 24148 28224 24200
rect 29644 24191 29696 24200
rect 27896 24080 27948 24089
rect 28356 24080 28408 24132
rect 29644 24157 29653 24191
rect 29653 24157 29687 24191
rect 29687 24157 29696 24191
rect 29644 24148 29696 24157
rect 31392 24191 31444 24200
rect 31392 24157 31401 24191
rect 31401 24157 31435 24191
rect 31435 24157 31444 24191
rect 31392 24148 31444 24157
rect 32864 24148 32916 24200
rect 33692 24191 33744 24200
rect 33692 24157 33701 24191
rect 33701 24157 33735 24191
rect 33735 24157 33744 24191
rect 33692 24148 33744 24157
rect 40132 24191 40184 24200
rect 40132 24157 40141 24191
rect 40141 24157 40175 24191
rect 40175 24157 40184 24191
rect 40132 24148 40184 24157
rect 30012 24123 30064 24132
rect 27160 24055 27212 24064
rect 27160 24021 27169 24055
rect 27169 24021 27203 24055
rect 27203 24021 27212 24055
rect 27160 24012 27212 24021
rect 29000 24055 29052 24064
rect 29000 24021 29009 24055
rect 29009 24021 29043 24055
rect 29043 24021 29052 24055
rect 30012 24089 30021 24123
rect 30021 24089 30055 24123
rect 30055 24089 30064 24123
rect 30012 24080 30064 24089
rect 40040 24080 40092 24132
rect 29000 24012 29052 24021
rect 33416 24012 33468 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 1584 23808 1636 23860
rect 12624 23808 12676 23860
rect 12900 23808 12952 23860
rect 13728 23808 13780 23860
rect 14280 23783 14332 23792
rect 2320 23536 2372 23588
rect 14280 23749 14289 23783
rect 14289 23749 14323 23783
rect 14323 23749 14332 23783
rect 14280 23740 14332 23749
rect 7380 23715 7432 23724
rect 7380 23681 7389 23715
rect 7389 23681 7423 23715
rect 7423 23681 7432 23715
rect 7380 23672 7432 23681
rect 9496 23672 9548 23724
rect 10416 23672 10468 23724
rect 11704 23715 11756 23724
rect 11704 23681 11713 23715
rect 11713 23681 11747 23715
rect 11747 23681 11756 23715
rect 11704 23672 11756 23681
rect 12532 23715 12584 23724
rect 12532 23681 12541 23715
rect 12541 23681 12575 23715
rect 12575 23681 12584 23715
rect 12532 23672 12584 23681
rect 12808 23715 12860 23724
rect 12808 23681 12817 23715
rect 12817 23681 12851 23715
rect 12851 23681 12860 23715
rect 12808 23672 12860 23681
rect 13360 23672 13412 23724
rect 14556 23715 14608 23724
rect 14556 23681 14565 23715
rect 14565 23681 14599 23715
rect 14599 23681 14608 23715
rect 17224 23740 17276 23792
rect 18512 23808 18564 23860
rect 20352 23851 20404 23860
rect 20352 23817 20361 23851
rect 20361 23817 20395 23851
rect 20395 23817 20404 23851
rect 20352 23808 20404 23817
rect 17960 23740 18012 23792
rect 19156 23740 19208 23792
rect 19432 23783 19484 23792
rect 19432 23749 19441 23783
rect 19441 23749 19475 23783
rect 19475 23749 19484 23783
rect 19432 23740 19484 23749
rect 20996 23808 21048 23860
rect 23296 23808 23348 23860
rect 25872 23808 25924 23860
rect 14556 23672 14608 23681
rect 17132 23715 17184 23724
rect 17132 23681 17141 23715
rect 17141 23681 17175 23715
rect 17175 23681 17184 23715
rect 17132 23672 17184 23681
rect 17500 23672 17552 23724
rect 18052 23672 18104 23724
rect 7564 23647 7616 23656
rect 7564 23613 7573 23647
rect 7573 23613 7607 23647
rect 7607 23613 7616 23647
rect 7564 23604 7616 23613
rect 9128 23647 9180 23656
rect 9128 23613 9137 23647
rect 9137 23613 9171 23647
rect 9171 23613 9180 23647
rect 9128 23604 9180 23613
rect 9588 23604 9640 23656
rect 11612 23647 11664 23656
rect 11612 23613 11621 23647
rect 11621 23613 11655 23647
rect 11655 23613 11664 23647
rect 11612 23604 11664 23613
rect 13544 23647 13596 23656
rect 13544 23613 13553 23647
rect 13553 23613 13587 23647
rect 13587 23613 13596 23647
rect 13544 23604 13596 23613
rect 2044 23511 2096 23520
rect 2044 23477 2053 23511
rect 2053 23477 2087 23511
rect 2087 23477 2096 23511
rect 2044 23468 2096 23477
rect 2688 23468 2740 23520
rect 11980 23536 12032 23588
rect 12624 23536 12676 23588
rect 17224 23604 17276 23656
rect 18328 23715 18380 23724
rect 18328 23681 18337 23715
rect 18337 23681 18371 23715
rect 18371 23681 18380 23715
rect 18512 23715 18564 23724
rect 18328 23672 18380 23681
rect 18512 23681 18521 23715
rect 18521 23681 18555 23715
rect 18555 23681 18564 23715
rect 18512 23672 18564 23681
rect 20076 23672 20128 23724
rect 23020 23740 23072 23792
rect 18420 23604 18472 23656
rect 20352 23604 20404 23656
rect 9864 23511 9916 23520
rect 9864 23477 9873 23511
rect 9873 23477 9907 23511
rect 9907 23477 9916 23511
rect 9864 23468 9916 23477
rect 12532 23511 12584 23520
rect 12532 23477 12541 23511
rect 12541 23477 12575 23511
rect 12575 23477 12584 23511
rect 12532 23468 12584 23477
rect 12716 23468 12768 23520
rect 14464 23511 14516 23520
rect 14464 23477 14473 23511
rect 14473 23477 14507 23511
rect 14507 23477 14516 23511
rect 14464 23468 14516 23477
rect 14740 23511 14792 23520
rect 14740 23477 14749 23511
rect 14749 23477 14783 23511
rect 14783 23477 14792 23511
rect 14740 23468 14792 23477
rect 16672 23511 16724 23520
rect 16672 23477 16681 23511
rect 16681 23477 16715 23511
rect 16715 23477 16724 23511
rect 16672 23468 16724 23477
rect 20628 23536 20680 23588
rect 20812 23715 20864 23724
rect 20812 23681 20826 23715
rect 20826 23681 20860 23715
rect 20860 23681 20864 23715
rect 20812 23672 20864 23681
rect 21180 23672 21232 23724
rect 23020 23604 23072 23656
rect 23848 23672 23900 23724
rect 23756 23604 23808 23656
rect 24400 23672 24452 23724
rect 25872 23672 25924 23724
rect 27896 23851 27948 23860
rect 27896 23817 27905 23851
rect 27905 23817 27939 23851
rect 27939 23817 27948 23851
rect 27896 23808 27948 23817
rect 28356 23808 28408 23860
rect 30012 23808 30064 23860
rect 30380 23808 30432 23860
rect 31576 23851 31628 23860
rect 31576 23817 31585 23851
rect 31585 23817 31619 23851
rect 31619 23817 31628 23851
rect 31576 23808 31628 23817
rect 32956 23808 33008 23860
rect 48044 23851 48096 23860
rect 48044 23817 48053 23851
rect 48053 23817 48087 23851
rect 48087 23817 48096 23851
rect 48044 23808 48096 23817
rect 26608 23740 26660 23792
rect 47308 23740 47360 23792
rect 47952 23783 48004 23792
rect 47952 23749 47961 23783
rect 47961 23749 47995 23783
rect 47995 23749 48004 23783
rect 47952 23740 48004 23749
rect 25780 23604 25832 23656
rect 26792 23672 26844 23724
rect 26976 23715 27028 23724
rect 26976 23681 26985 23715
rect 26985 23681 27019 23715
rect 27019 23681 27028 23715
rect 26976 23672 27028 23681
rect 27160 23715 27212 23724
rect 27160 23681 27169 23715
rect 27169 23681 27203 23715
rect 27203 23681 27212 23715
rect 27160 23672 27212 23681
rect 27804 23672 27856 23724
rect 28080 23604 28132 23656
rect 28356 23715 28408 23724
rect 28356 23681 28365 23715
rect 28365 23681 28399 23715
rect 28399 23681 28408 23715
rect 28356 23672 28408 23681
rect 29368 23715 29420 23724
rect 21916 23536 21968 23588
rect 22928 23579 22980 23588
rect 22928 23545 22937 23579
rect 22937 23545 22971 23579
rect 22971 23545 22980 23579
rect 22928 23536 22980 23545
rect 24676 23536 24728 23588
rect 26792 23536 26844 23588
rect 29368 23681 29377 23715
rect 29377 23681 29411 23715
rect 29411 23681 29420 23715
rect 29368 23672 29420 23681
rect 30288 23672 30340 23724
rect 30472 23715 30524 23724
rect 30472 23681 30506 23715
rect 30506 23681 30524 23715
rect 30472 23672 30524 23681
rect 32496 23672 32548 23724
rect 30196 23647 30248 23656
rect 30196 23613 30205 23647
rect 30205 23613 30239 23647
rect 30239 23613 30248 23647
rect 30196 23604 30248 23613
rect 33232 23647 33284 23656
rect 33232 23613 33241 23647
rect 33241 23613 33275 23647
rect 33275 23613 33284 23647
rect 33232 23604 33284 23613
rect 33416 23647 33468 23656
rect 33416 23613 33425 23647
rect 33425 23613 33459 23647
rect 33459 23613 33468 23647
rect 33416 23604 33468 23613
rect 33784 23647 33836 23656
rect 33784 23613 33793 23647
rect 33793 23613 33827 23647
rect 33827 23613 33836 23647
rect 33784 23604 33836 23613
rect 28908 23536 28960 23588
rect 17684 23468 17736 23520
rect 17868 23511 17920 23520
rect 17868 23477 17877 23511
rect 17877 23477 17911 23511
rect 17911 23477 17920 23511
rect 17868 23468 17920 23477
rect 19432 23468 19484 23520
rect 21548 23468 21600 23520
rect 23664 23468 23716 23520
rect 26240 23468 26292 23520
rect 29552 23468 29604 23520
rect 30380 23468 30432 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 7564 23264 7616 23316
rect 9496 23307 9548 23316
rect 9496 23273 9505 23307
rect 9505 23273 9539 23307
rect 9539 23273 9548 23307
rect 9496 23264 9548 23273
rect 9680 23307 9732 23316
rect 9680 23273 9689 23307
rect 9689 23273 9723 23307
rect 9723 23273 9732 23307
rect 9680 23264 9732 23273
rect 9772 23264 9824 23316
rect 2504 23196 2556 23248
rect 4712 23196 4764 23248
rect 2044 23128 2096 23180
rect 2780 23171 2832 23180
rect 2780 23137 2789 23171
rect 2789 23137 2823 23171
rect 2823 23137 2832 23171
rect 2780 23128 2832 23137
rect 2596 22992 2648 23044
rect 10324 23196 10376 23248
rect 11612 23264 11664 23316
rect 12532 23307 12584 23316
rect 12532 23273 12541 23307
rect 12541 23273 12575 23307
rect 12575 23273 12584 23307
rect 12532 23264 12584 23273
rect 12992 23307 13044 23316
rect 12992 23273 13001 23307
rect 13001 23273 13035 23307
rect 13035 23273 13044 23307
rect 12992 23264 13044 23273
rect 14280 23307 14332 23316
rect 14280 23273 14289 23307
rect 14289 23273 14323 23307
rect 14323 23273 14332 23307
rect 14280 23264 14332 23273
rect 14464 23307 14516 23316
rect 14464 23273 14473 23307
rect 14473 23273 14507 23307
rect 14507 23273 14516 23307
rect 14464 23264 14516 23273
rect 16580 23196 16632 23248
rect 18328 23196 18380 23248
rect 20812 23196 20864 23248
rect 23940 23264 23992 23316
rect 24308 23264 24360 23316
rect 25688 23264 25740 23316
rect 25964 23264 26016 23316
rect 28356 23264 28408 23316
rect 30472 23264 30524 23316
rect 10416 23171 10468 23180
rect 7748 23103 7800 23112
rect 7748 23069 7757 23103
rect 7757 23069 7791 23103
rect 7791 23069 7800 23103
rect 7748 23060 7800 23069
rect 8024 23060 8076 23112
rect 10416 23137 10425 23171
rect 10425 23137 10459 23171
rect 10459 23137 10468 23171
rect 10416 23128 10468 23137
rect 12624 23171 12676 23180
rect 12624 23137 12633 23171
rect 12633 23137 12667 23171
rect 12667 23137 12676 23171
rect 12624 23128 12676 23137
rect 10324 23103 10376 23112
rect 10324 23069 10333 23103
rect 10333 23069 10367 23103
rect 10367 23069 10376 23103
rect 10324 23060 10376 23069
rect 14740 23128 14792 23180
rect 13084 23060 13136 23112
rect 15568 23103 15620 23112
rect 9588 22992 9640 23044
rect 14096 23035 14148 23044
rect 14096 23001 14131 23035
rect 14131 23001 14148 23035
rect 14096 22992 14148 23001
rect 9772 22924 9824 22976
rect 13636 22924 13688 22976
rect 14372 22992 14424 23044
rect 15568 23069 15577 23103
rect 15577 23069 15611 23103
rect 15611 23069 15620 23103
rect 15568 23060 15620 23069
rect 16672 23060 16724 23112
rect 18788 23060 18840 23112
rect 19156 23060 19208 23112
rect 17960 22992 18012 23044
rect 18052 22992 18104 23044
rect 22928 23060 22980 23112
rect 23296 23060 23348 23112
rect 24032 23128 24084 23180
rect 24492 23171 24544 23180
rect 24492 23137 24501 23171
rect 24501 23137 24535 23171
rect 24535 23137 24544 23171
rect 24492 23128 24544 23137
rect 24584 23060 24636 23112
rect 14464 22924 14516 22976
rect 20720 22992 20772 23044
rect 20812 22992 20864 23044
rect 21732 22992 21784 23044
rect 24400 23035 24452 23044
rect 24400 23001 24409 23035
rect 24409 23001 24443 23035
rect 24443 23001 24452 23035
rect 24400 22992 24452 23001
rect 28080 23196 28132 23248
rect 28908 23128 28960 23180
rect 29092 23128 29144 23180
rect 29000 23060 29052 23112
rect 29828 23060 29880 23112
rect 30380 23103 30432 23112
rect 30380 23069 30389 23103
rect 30389 23069 30423 23103
rect 30423 23069 30432 23103
rect 30380 23060 30432 23069
rect 30656 23060 30708 23112
rect 32496 23060 32548 23112
rect 21180 22967 21232 22976
rect 21180 22933 21189 22967
rect 21189 22933 21223 22967
rect 21223 22933 21232 22967
rect 21180 22924 21232 22933
rect 23572 22924 23624 22976
rect 24216 22924 24268 22976
rect 26240 22924 26292 22976
rect 26976 22992 27028 23044
rect 27252 22992 27304 23044
rect 29368 22992 29420 23044
rect 30932 22924 30984 22976
rect 31116 22967 31168 22976
rect 31116 22933 31125 22967
rect 31125 22933 31159 22967
rect 31159 22933 31168 22967
rect 31116 22924 31168 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 2596 22763 2648 22772
rect 2596 22729 2605 22763
rect 2605 22729 2639 22763
rect 2639 22729 2648 22763
rect 2596 22720 2648 22729
rect 1492 22652 1544 22704
rect 12808 22695 12860 22704
rect 12808 22661 12817 22695
rect 12817 22661 12851 22695
rect 12851 22661 12860 22695
rect 12808 22652 12860 22661
rect 13636 22695 13688 22704
rect 13636 22661 13645 22695
rect 13645 22661 13679 22695
rect 13679 22661 13688 22695
rect 13636 22652 13688 22661
rect 14280 22695 14332 22704
rect 14280 22661 14289 22695
rect 14289 22661 14323 22695
rect 14323 22661 14332 22695
rect 14280 22652 14332 22661
rect 14464 22652 14516 22704
rect 17224 22652 17276 22704
rect 17868 22652 17920 22704
rect 1860 22627 1912 22636
rect 1860 22593 1869 22627
rect 1869 22593 1903 22627
rect 1903 22593 1912 22627
rect 1860 22584 1912 22593
rect 2504 22627 2556 22636
rect 2504 22593 2513 22627
rect 2513 22593 2547 22627
rect 2547 22593 2556 22627
rect 2504 22584 2556 22593
rect 1952 22516 2004 22568
rect 2596 22516 2648 22568
rect 13268 22584 13320 22636
rect 13360 22627 13412 22636
rect 13360 22593 13369 22627
rect 13369 22593 13403 22627
rect 13403 22593 13412 22627
rect 14096 22627 14148 22636
rect 13360 22584 13412 22593
rect 14096 22593 14105 22627
rect 14105 22593 14139 22627
rect 14139 22593 14148 22627
rect 14096 22584 14148 22593
rect 13176 22516 13228 22568
rect 13452 22559 13504 22568
rect 13452 22525 13461 22559
rect 13461 22525 13495 22559
rect 13495 22525 13504 22559
rect 13452 22516 13504 22525
rect 13636 22559 13688 22568
rect 13636 22525 13645 22559
rect 13645 22525 13679 22559
rect 13679 22525 13688 22559
rect 13636 22516 13688 22525
rect 14372 22627 14424 22636
rect 14372 22593 14381 22627
rect 14381 22593 14415 22627
rect 14415 22593 14424 22627
rect 14372 22584 14424 22593
rect 21180 22652 21232 22704
rect 23848 22695 23900 22704
rect 23848 22661 23857 22695
rect 23857 22661 23891 22695
rect 23891 22661 23900 22695
rect 23848 22652 23900 22661
rect 24676 22652 24728 22704
rect 19156 22584 19208 22636
rect 21824 22627 21876 22636
rect 15568 22516 15620 22568
rect 19248 22559 19300 22568
rect 14556 22448 14608 22500
rect 1952 22423 2004 22432
rect 1952 22389 1961 22423
rect 1961 22389 1995 22423
rect 1995 22389 2004 22423
rect 1952 22380 2004 22389
rect 19248 22525 19257 22559
rect 19257 22525 19291 22559
rect 19291 22525 19300 22559
rect 19248 22516 19300 22525
rect 18788 22491 18840 22500
rect 18788 22457 18797 22491
rect 18797 22457 18831 22491
rect 18831 22457 18840 22491
rect 18788 22448 18840 22457
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 22100 22627 22152 22636
rect 22100 22593 22134 22627
rect 22134 22593 22152 22627
rect 22100 22584 22152 22593
rect 23020 22584 23072 22636
rect 24584 22584 24636 22636
rect 24860 22627 24912 22636
rect 24860 22593 24869 22627
rect 24869 22593 24903 22627
rect 24903 22593 24912 22627
rect 24860 22584 24912 22593
rect 25136 22627 25188 22636
rect 25136 22593 25145 22627
rect 25145 22593 25179 22627
rect 25179 22593 25188 22627
rect 25136 22584 25188 22593
rect 26240 22652 26292 22704
rect 26884 22652 26936 22704
rect 27252 22627 27304 22636
rect 27252 22593 27261 22627
rect 27261 22593 27295 22627
rect 27295 22593 27304 22627
rect 27252 22584 27304 22593
rect 29460 22627 29512 22636
rect 29460 22593 29469 22627
rect 29469 22593 29503 22627
rect 29503 22593 29512 22627
rect 29460 22584 29512 22593
rect 30564 22720 30616 22772
rect 30840 22720 30892 22772
rect 29828 22652 29880 22704
rect 29736 22627 29788 22636
rect 29736 22593 29745 22627
rect 29745 22593 29779 22627
rect 29779 22593 29788 22627
rect 29736 22584 29788 22593
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 46940 22652 46992 22704
rect 25320 22516 25372 22568
rect 34244 22627 34296 22636
rect 34244 22593 34253 22627
rect 34253 22593 34287 22627
rect 34287 22593 34296 22627
rect 34244 22584 34296 22593
rect 48136 22627 48188 22636
rect 48136 22593 48145 22627
rect 48145 22593 48179 22627
rect 48179 22593 48188 22627
rect 48136 22584 48188 22593
rect 21364 22448 21416 22500
rect 18696 22380 18748 22432
rect 21732 22380 21784 22432
rect 23940 22448 23992 22500
rect 25228 22380 25280 22432
rect 25780 22380 25832 22432
rect 29460 22380 29512 22432
rect 33876 22380 33928 22432
rect 34152 22448 34204 22500
rect 34520 22380 34572 22432
rect 47584 22380 47636 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 1952 22176 2004 22228
rect 13360 22176 13412 22228
rect 14280 22219 14332 22228
rect 14280 22185 14289 22219
rect 14289 22185 14323 22219
rect 14323 22185 14332 22219
rect 14280 22176 14332 22185
rect 14464 22151 14516 22160
rect 14464 22117 14473 22151
rect 14473 22117 14507 22151
rect 14507 22117 14516 22151
rect 20720 22176 20772 22228
rect 21824 22176 21876 22228
rect 23756 22176 23808 22228
rect 24400 22219 24452 22228
rect 24400 22185 24409 22219
rect 24409 22185 24443 22219
rect 24443 22185 24452 22219
rect 24400 22176 24452 22185
rect 25136 22176 25188 22228
rect 14464 22108 14516 22117
rect 22284 22108 22336 22160
rect 1676 22040 1728 22092
rect 18052 22040 18104 22092
rect 7012 21972 7064 22024
rect 8208 21972 8260 22024
rect 10232 22015 10284 22024
rect 10232 21981 10241 22015
rect 10241 21981 10275 22015
rect 10275 21981 10284 22015
rect 10232 21972 10284 21981
rect 12992 21972 13044 22024
rect 14188 21972 14240 22024
rect 14372 21972 14424 22024
rect 9220 21904 9272 21956
rect 11612 21904 11664 21956
rect 9772 21836 9824 21888
rect 10600 21836 10652 21888
rect 11244 21836 11296 21888
rect 13084 21904 13136 21956
rect 18420 22015 18472 22024
rect 18420 21981 18429 22015
rect 18429 21981 18463 22015
rect 18463 21981 18472 22015
rect 18420 21972 18472 21981
rect 18512 22015 18564 22024
rect 18512 21981 18521 22015
rect 18521 21981 18555 22015
rect 18555 21981 18564 22015
rect 18512 21972 18564 21981
rect 18788 21972 18840 22024
rect 18880 21972 18932 22024
rect 20720 21972 20772 22024
rect 20996 21972 21048 22024
rect 21916 22040 21968 22092
rect 21732 21972 21784 22024
rect 22652 21972 22704 22024
rect 24492 22108 24544 22160
rect 23848 22015 23900 22024
rect 23848 21981 23857 22015
rect 23857 21981 23891 22015
rect 23891 21981 23900 22015
rect 23848 21972 23900 21981
rect 20260 21904 20312 21956
rect 23756 21904 23808 21956
rect 25504 22176 25556 22228
rect 29736 22176 29788 22228
rect 34152 22176 34204 22228
rect 34612 22176 34664 22228
rect 29092 22108 29144 22160
rect 30656 22108 30708 22160
rect 32036 22108 32088 22160
rect 31116 22040 31168 22092
rect 34244 22108 34296 22160
rect 36636 22176 36688 22228
rect 47768 22176 47820 22228
rect 47400 22083 47452 22092
rect 24400 21947 24452 21956
rect 24400 21913 24409 21947
rect 24409 21913 24443 21947
rect 24443 21913 24452 21947
rect 24400 21904 24452 21913
rect 25228 21972 25280 22024
rect 25596 22015 25648 22024
rect 25596 21981 25605 22015
rect 25605 21981 25639 22015
rect 25639 21981 25648 22015
rect 27620 22015 27672 22024
rect 25596 21972 25648 21981
rect 27620 21981 27629 22015
rect 27629 21981 27663 22015
rect 27663 21981 27672 22015
rect 27620 21972 27672 21981
rect 29552 22015 29604 22024
rect 29552 21981 29561 22015
rect 29561 21981 29595 22015
rect 29595 21981 29604 22015
rect 29552 21972 29604 21981
rect 47400 22049 47409 22083
rect 47409 22049 47443 22083
rect 47443 22049 47452 22083
rect 47400 22040 47452 22049
rect 13452 21836 13504 21888
rect 13636 21836 13688 21888
rect 14372 21836 14424 21888
rect 15844 21836 15896 21888
rect 20628 21879 20680 21888
rect 20628 21845 20637 21879
rect 20637 21845 20671 21879
rect 20671 21845 20680 21879
rect 20628 21836 20680 21845
rect 24584 21836 24636 21888
rect 25412 21904 25464 21956
rect 27160 21836 27212 21888
rect 28264 21904 28316 21956
rect 29920 21904 29972 21956
rect 31300 21904 31352 21956
rect 32680 21947 32732 21956
rect 32680 21913 32689 21947
rect 32689 21913 32723 21947
rect 32723 21913 32732 21947
rect 32680 21904 32732 21913
rect 32864 21947 32916 21956
rect 32864 21913 32873 21947
rect 32873 21913 32907 21947
rect 32907 21913 32916 21947
rect 32864 21904 32916 21913
rect 33968 22015 34020 22024
rect 33968 21981 33977 22015
rect 33977 21981 34011 22015
rect 34011 21981 34020 22015
rect 33968 21972 34020 21981
rect 34152 22015 34204 22024
rect 34152 21981 34161 22015
rect 34161 21981 34195 22015
rect 34195 21981 34204 22015
rect 34704 22015 34756 22024
rect 34152 21972 34204 21981
rect 34704 21981 34713 22015
rect 34713 21981 34747 22015
rect 34747 21981 34756 22015
rect 34704 21972 34756 21981
rect 47584 21972 47636 22024
rect 47860 22015 47912 22024
rect 47860 21981 47869 22015
rect 47869 21981 47903 22015
rect 47903 21981 47912 22015
rect 47860 21972 47912 21981
rect 34520 21904 34572 21956
rect 29552 21836 29604 21888
rect 36084 21879 36136 21888
rect 36084 21845 36093 21879
rect 36093 21845 36127 21879
rect 36127 21845 36136 21879
rect 36084 21836 36136 21845
rect 36544 21836 36596 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 8208 21632 8260 21684
rect 11612 21675 11664 21684
rect 11612 21641 11621 21675
rect 11621 21641 11655 21675
rect 11655 21641 11664 21675
rect 11612 21632 11664 21641
rect 13728 21632 13780 21684
rect 18512 21632 18564 21684
rect 9404 21564 9456 21616
rect 2412 21496 2464 21548
rect 9496 21496 9548 21548
rect 9772 21539 9824 21548
rect 9772 21505 9781 21539
rect 9781 21505 9815 21539
rect 9815 21505 9824 21539
rect 9772 21496 9824 21505
rect 7472 21471 7524 21480
rect 7472 21437 7481 21471
rect 7481 21437 7515 21471
rect 7515 21437 7524 21471
rect 7472 21428 7524 21437
rect 10232 21496 10284 21548
rect 12992 21539 13044 21548
rect 12992 21505 13001 21539
rect 13001 21505 13035 21539
rect 13035 21505 13044 21539
rect 12992 21496 13044 21505
rect 13360 21496 13412 21548
rect 9496 21360 9548 21412
rect 14280 21471 14332 21480
rect 14280 21437 14289 21471
rect 14289 21437 14323 21471
rect 14323 21437 14332 21471
rect 14280 21428 14332 21437
rect 20628 21564 20680 21616
rect 20812 21564 20864 21616
rect 17868 21539 17920 21548
rect 17868 21505 17877 21539
rect 17877 21505 17911 21539
rect 17911 21505 17920 21539
rect 17868 21496 17920 21505
rect 19248 21496 19300 21548
rect 19432 21496 19484 21548
rect 20076 21496 20128 21548
rect 26240 21632 26292 21684
rect 28264 21675 28316 21684
rect 20996 21564 21048 21616
rect 21548 21496 21600 21548
rect 23664 21496 23716 21548
rect 24124 21496 24176 21548
rect 25780 21539 25832 21548
rect 25780 21505 25789 21539
rect 25789 21505 25823 21539
rect 25823 21505 25832 21539
rect 25780 21496 25832 21505
rect 26148 21564 26200 21616
rect 26976 21607 27028 21616
rect 26976 21573 26985 21607
rect 26985 21573 27019 21607
rect 27019 21573 27028 21607
rect 26976 21564 27028 21573
rect 27160 21539 27212 21548
rect 21180 21428 21232 21480
rect 21824 21428 21876 21480
rect 24032 21428 24084 21480
rect 24768 21428 24820 21480
rect 25412 21471 25464 21480
rect 25412 21437 25421 21471
rect 25421 21437 25455 21471
rect 25455 21437 25464 21471
rect 25412 21428 25464 21437
rect 27160 21505 27169 21539
rect 27169 21505 27203 21539
rect 27203 21505 27212 21539
rect 27160 21496 27212 21505
rect 28264 21641 28273 21675
rect 28273 21641 28307 21675
rect 28307 21641 28316 21675
rect 28264 21632 28316 21641
rect 30564 21675 30616 21684
rect 30564 21641 30573 21675
rect 30573 21641 30607 21675
rect 30607 21641 30616 21675
rect 30564 21632 30616 21641
rect 29184 21564 29236 21616
rect 29368 21607 29420 21616
rect 29368 21573 29377 21607
rect 29377 21573 29411 21607
rect 29411 21573 29420 21607
rect 29368 21564 29420 21573
rect 29552 21607 29604 21616
rect 29552 21573 29561 21607
rect 29561 21573 29595 21607
rect 29595 21573 29604 21607
rect 29552 21564 29604 21573
rect 29644 21564 29696 21616
rect 47768 21632 47820 21684
rect 28908 21539 28960 21548
rect 28080 21428 28132 21480
rect 28908 21505 28917 21539
rect 28917 21505 28951 21539
rect 28951 21505 28960 21539
rect 28908 21496 28960 21505
rect 30840 21496 30892 21548
rect 34704 21564 34756 21616
rect 47952 21607 48004 21616
rect 47952 21573 47961 21607
rect 47961 21573 47995 21607
rect 47995 21573 48004 21607
rect 47952 21564 48004 21573
rect 33876 21496 33928 21548
rect 15660 21360 15712 21412
rect 17316 21403 17368 21412
rect 17316 21369 17325 21403
rect 17325 21369 17359 21403
rect 17359 21369 17368 21403
rect 17316 21360 17368 21369
rect 18420 21360 18472 21412
rect 19248 21360 19300 21412
rect 24584 21360 24636 21412
rect 29644 21360 29696 21412
rect 13084 21292 13136 21344
rect 13452 21292 13504 21344
rect 14004 21292 14056 21344
rect 17500 21292 17552 21344
rect 19432 21292 19484 21344
rect 23480 21335 23532 21344
rect 23480 21301 23489 21335
rect 23489 21301 23523 21335
rect 23523 21301 23532 21335
rect 23480 21292 23532 21301
rect 24492 21292 24544 21344
rect 32680 21428 32732 21480
rect 31852 21292 31904 21344
rect 32864 21292 32916 21344
rect 48044 21335 48096 21344
rect 48044 21301 48053 21335
rect 48053 21301 48087 21335
rect 48087 21301 48096 21335
rect 48044 21292 48096 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4620 21088 4672 21140
rect 3976 21020 4028 21072
rect 15660 21063 15712 21072
rect 4068 20952 4120 21004
rect 10600 20995 10652 21004
rect 10600 20961 10609 20995
rect 10609 20961 10643 20995
rect 10643 20961 10652 20995
rect 10600 20952 10652 20961
rect 15660 21029 15669 21063
rect 15669 21029 15703 21063
rect 15703 21029 15712 21063
rect 15660 21020 15712 21029
rect 9036 20884 9088 20936
rect 9309 20924 9361 20933
rect 9309 20890 9318 20924
rect 9318 20890 9352 20924
rect 9352 20890 9361 20924
rect 9309 20881 9361 20890
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 6460 20859 6512 20868
rect 6460 20825 6469 20859
rect 6469 20825 6503 20859
rect 6503 20825 6512 20859
rect 6460 20816 6512 20825
rect 13176 20884 13228 20936
rect 10784 20816 10836 20868
rect 14556 20859 14608 20868
rect 14556 20825 14590 20859
rect 14590 20825 14608 20859
rect 14556 20816 14608 20825
rect 8208 20748 8260 20800
rect 8944 20791 8996 20800
rect 8944 20757 8953 20791
rect 8953 20757 8987 20791
rect 8987 20757 8996 20791
rect 8944 20748 8996 20757
rect 9496 20748 9548 20800
rect 16488 20816 16540 20868
rect 18696 21088 18748 21140
rect 20996 21088 21048 21140
rect 21548 21020 21600 21072
rect 17868 20952 17920 21004
rect 21456 20952 21508 21004
rect 25136 21088 25188 21140
rect 33968 21131 34020 21140
rect 29460 21020 29512 21072
rect 31116 21020 31168 21072
rect 33968 21097 33977 21131
rect 33977 21097 34011 21131
rect 34011 21097 34020 21131
rect 33968 21088 34020 21097
rect 20720 20927 20772 20936
rect 20720 20893 20729 20927
rect 20729 20893 20763 20927
rect 20763 20893 20772 20927
rect 20720 20884 20772 20893
rect 27160 20952 27212 21004
rect 36544 21020 36596 21072
rect 22100 20884 22152 20936
rect 23480 20884 23532 20936
rect 16764 20748 16816 20800
rect 16856 20748 16908 20800
rect 18788 20748 18840 20800
rect 20996 20748 21048 20800
rect 21456 20748 21508 20800
rect 22652 20791 22704 20800
rect 22652 20757 22661 20791
rect 22661 20757 22695 20791
rect 22695 20757 22704 20791
rect 22652 20748 22704 20757
rect 24032 20816 24084 20868
rect 24492 20884 24544 20936
rect 26240 20927 26292 20936
rect 26240 20893 26249 20927
rect 26249 20893 26283 20927
rect 26283 20893 26292 20927
rect 26240 20884 26292 20893
rect 31208 20884 31260 20936
rect 26148 20816 26200 20868
rect 28724 20859 28776 20868
rect 28724 20825 28733 20859
rect 28733 20825 28767 20859
rect 28767 20825 28776 20859
rect 28724 20816 28776 20825
rect 30656 20816 30708 20868
rect 32036 20884 32088 20936
rect 32588 20927 32640 20936
rect 32588 20893 32597 20927
rect 32597 20893 32631 20927
rect 32631 20893 32640 20927
rect 32588 20884 32640 20893
rect 32680 20884 32732 20936
rect 33692 20884 33744 20936
rect 36084 20884 36136 20936
rect 27988 20748 28040 20800
rect 32128 20748 32180 20800
rect 32312 20816 32364 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 6460 20587 6512 20596
rect 6460 20553 6469 20587
rect 6469 20553 6503 20587
rect 6503 20553 6512 20587
rect 6460 20544 6512 20553
rect 8208 20544 8260 20596
rect 6368 20451 6420 20460
rect 6368 20417 6377 20451
rect 6377 20417 6411 20451
rect 6411 20417 6420 20451
rect 6368 20408 6420 20417
rect 7472 20476 7524 20528
rect 7840 20476 7892 20528
rect 9404 20544 9456 20596
rect 14556 20544 14608 20596
rect 16764 20544 16816 20596
rect 23480 20544 23532 20596
rect 8944 20408 8996 20460
rect 9220 20451 9272 20460
rect 9220 20417 9229 20451
rect 9229 20417 9263 20451
rect 9263 20417 9272 20451
rect 9220 20408 9272 20417
rect 10600 20451 10652 20460
rect 10600 20417 10609 20451
rect 10609 20417 10643 20451
rect 10643 20417 10652 20451
rect 10600 20408 10652 20417
rect 10784 20451 10836 20460
rect 10784 20417 10793 20451
rect 10793 20417 10827 20451
rect 10827 20417 10836 20451
rect 10784 20408 10836 20417
rect 10968 20451 11020 20460
rect 10968 20417 10977 20451
rect 10977 20417 11011 20451
rect 11011 20417 11020 20451
rect 10968 20408 11020 20417
rect 11980 20408 12032 20460
rect 12348 20451 12400 20460
rect 12348 20417 12357 20451
rect 12357 20417 12391 20451
rect 12391 20417 12400 20451
rect 12348 20408 12400 20417
rect 12440 20451 12492 20460
rect 12440 20417 12449 20451
rect 12449 20417 12483 20451
rect 12483 20417 12492 20451
rect 12624 20451 12676 20460
rect 12440 20408 12492 20417
rect 12624 20417 12633 20451
rect 12633 20417 12667 20451
rect 12667 20417 12676 20451
rect 12624 20408 12676 20417
rect 12072 20340 12124 20392
rect 6368 20204 6420 20256
rect 12256 20272 12308 20324
rect 13820 20451 13872 20460
rect 13820 20417 13829 20451
rect 13829 20417 13863 20451
rect 13863 20417 13872 20451
rect 13820 20408 13872 20417
rect 14004 20451 14056 20460
rect 14004 20417 14013 20451
rect 14013 20417 14047 20451
rect 14047 20417 14056 20451
rect 14004 20408 14056 20417
rect 13912 20272 13964 20324
rect 14924 20451 14976 20460
rect 14924 20417 14933 20451
rect 14933 20417 14967 20451
rect 14967 20417 14976 20451
rect 14924 20408 14976 20417
rect 15108 20451 15160 20460
rect 15108 20417 15117 20451
rect 15117 20417 15151 20451
rect 15151 20417 15160 20451
rect 15108 20408 15160 20417
rect 15844 20451 15896 20460
rect 15844 20417 15853 20451
rect 15853 20417 15887 20451
rect 15887 20417 15896 20451
rect 15844 20408 15896 20417
rect 16764 20408 16816 20460
rect 17684 20476 17736 20528
rect 20260 20476 20312 20528
rect 27988 20519 28040 20528
rect 15936 20340 15988 20392
rect 11152 20204 11204 20256
rect 13452 20204 13504 20256
rect 17316 20451 17368 20460
rect 17316 20417 17325 20451
rect 17325 20417 17359 20451
rect 17359 20417 17368 20451
rect 18052 20451 18104 20460
rect 17316 20408 17368 20417
rect 18052 20417 18061 20451
rect 18061 20417 18095 20451
rect 18095 20417 18104 20451
rect 18052 20408 18104 20417
rect 20076 20408 20128 20460
rect 27988 20485 27997 20519
rect 27997 20485 28031 20519
rect 28031 20485 28040 20519
rect 27988 20476 28040 20485
rect 29276 20476 29328 20528
rect 29736 20476 29788 20528
rect 31668 20476 31720 20528
rect 18328 20340 18380 20392
rect 19248 20340 19300 20392
rect 20720 20451 20772 20460
rect 20720 20417 20729 20451
rect 20729 20417 20763 20451
rect 20763 20417 20772 20451
rect 20720 20408 20772 20417
rect 20996 20408 21048 20460
rect 22100 20408 22152 20460
rect 23296 20451 23348 20460
rect 23296 20417 23305 20451
rect 23305 20417 23339 20451
rect 23339 20417 23348 20451
rect 23296 20408 23348 20417
rect 23480 20408 23532 20460
rect 30196 20451 30248 20460
rect 21732 20340 21784 20392
rect 23940 20340 23992 20392
rect 17500 20272 17552 20324
rect 26608 20272 26660 20324
rect 17684 20247 17736 20256
rect 17684 20213 17693 20247
rect 17693 20213 17727 20247
rect 17727 20213 17736 20247
rect 17684 20204 17736 20213
rect 18512 20204 18564 20256
rect 18604 20204 18656 20256
rect 19892 20204 19944 20256
rect 21456 20204 21508 20256
rect 21916 20204 21968 20256
rect 22652 20204 22704 20256
rect 23204 20204 23256 20256
rect 24032 20204 24084 20256
rect 24308 20204 24360 20256
rect 30196 20417 30205 20451
rect 30205 20417 30239 20451
rect 30239 20417 30248 20451
rect 30196 20408 30248 20417
rect 30288 20408 30340 20460
rect 34704 20476 34756 20528
rect 48044 20476 48096 20528
rect 32220 20408 32272 20460
rect 32680 20408 32732 20460
rect 34244 20451 34296 20460
rect 34244 20417 34253 20451
rect 34253 20417 34287 20451
rect 34287 20417 34296 20451
rect 34244 20408 34296 20417
rect 34428 20451 34480 20460
rect 34428 20417 34437 20451
rect 34437 20417 34471 20451
rect 34471 20417 34480 20451
rect 34428 20408 34480 20417
rect 34612 20451 34664 20460
rect 34612 20417 34621 20451
rect 34621 20417 34655 20451
rect 34655 20417 34664 20451
rect 34612 20408 34664 20417
rect 31392 20272 31444 20324
rect 34520 20340 34572 20392
rect 41604 20272 41656 20324
rect 33968 20247 34020 20256
rect 33968 20213 33977 20247
rect 33977 20213 34011 20247
rect 34011 20213 34020 20247
rect 33968 20204 34020 20213
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 10784 20000 10836 20052
rect 13820 20000 13872 20052
rect 14924 20000 14976 20052
rect 12256 19932 12308 19984
rect 17684 20000 17736 20052
rect 47032 20000 47084 20052
rect 12072 19864 12124 19916
rect 12348 19864 12400 19916
rect 16120 19864 16172 19916
rect 20260 19932 20312 19984
rect 20536 19932 20588 19984
rect 25780 19975 25832 19984
rect 25780 19941 25789 19975
rect 25789 19941 25823 19975
rect 25823 19941 25832 19975
rect 25780 19932 25832 19941
rect 26792 19932 26844 19984
rect 31208 19932 31260 19984
rect 1860 19796 1912 19848
rect 7840 19728 7892 19780
rect 11152 19796 11204 19848
rect 11796 19796 11848 19848
rect 12992 19796 13044 19848
rect 14280 19839 14332 19848
rect 10600 19728 10652 19780
rect 13360 19771 13412 19780
rect 13360 19737 13369 19771
rect 13369 19737 13403 19771
rect 13403 19737 13412 19771
rect 13360 19728 13412 19737
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 16856 19796 16908 19848
rect 15936 19728 15988 19780
rect 17684 19796 17736 19848
rect 18236 19796 18288 19848
rect 18512 19839 18564 19848
rect 18512 19805 18521 19839
rect 18521 19805 18555 19839
rect 18555 19805 18564 19839
rect 18512 19796 18564 19805
rect 18696 19839 18748 19848
rect 18696 19805 18705 19839
rect 18705 19805 18739 19839
rect 18739 19805 18748 19839
rect 19248 19839 19300 19848
rect 18696 19796 18748 19805
rect 19248 19805 19257 19839
rect 19257 19805 19291 19839
rect 19291 19805 19300 19839
rect 19248 19796 19300 19805
rect 26608 19864 26660 19916
rect 17500 19728 17552 19780
rect 4068 19660 4120 19712
rect 8208 19660 8260 19712
rect 10416 19660 10468 19712
rect 12808 19660 12860 19712
rect 16856 19660 16908 19712
rect 19892 19796 19944 19848
rect 20260 19796 20312 19848
rect 21180 19839 21232 19848
rect 21180 19805 21189 19839
rect 21189 19805 21223 19839
rect 21223 19805 21232 19839
rect 21180 19796 21232 19805
rect 21456 19839 21508 19848
rect 21456 19805 21490 19839
rect 21490 19805 21508 19839
rect 21456 19796 21508 19805
rect 25596 19796 25648 19848
rect 27620 19796 27672 19848
rect 31392 19864 31444 19916
rect 30748 19796 30800 19848
rect 34428 19932 34480 19984
rect 34704 19907 34756 19916
rect 34704 19873 34713 19907
rect 34713 19873 34747 19907
rect 34747 19873 34756 19907
rect 34704 19864 34756 19873
rect 47768 19864 47820 19916
rect 22560 19703 22612 19712
rect 22560 19669 22569 19703
rect 22569 19669 22603 19703
rect 22603 19669 22612 19703
rect 22560 19660 22612 19669
rect 22652 19660 22704 19712
rect 23664 19660 23716 19712
rect 26056 19728 26108 19780
rect 27804 19771 27856 19780
rect 24768 19660 24820 19712
rect 27804 19737 27813 19771
rect 27813 19737 27847 19771
rect 27847 19737 27856 19771
rect 27804 19728 27856 19737
rect 28632 19728 28684 19780
rect 26792 19660 26844 19712
rect 32312 19796 32364 19848
rect 33232 19796 33284 19848
rect 33692 19839 33744 19848
rect 33692 19805 33701 19839
rect 33701 19805 33735 19839
rect 33735 19805 33744 19839
rect 33692 19796 33744 19805
rect 33876 19839 33928 19848
rect 33876 19805 33885 19839
rect 33885 19805 33919 19839
rect 33919 19805 33928 19839
rect 33876 19796 33928 19805
rect 33968 19796 34020 19848
rect 46756 19728 46808 19780
rect 48136 19771 48188 19780
rect 48136 19737 48145 19771
rect 48145 19737 48179 19771
rect 48179 19737 48188 19771
rect 48136 19728 48188 19737
rect 30012 19660 30064 19712
rect 31760 19703 31812 19712
rect 31760 19669 31769 19703
rect 31769 19669 31803 19703
rect 31803 19669 31812 19703
rect 31760 19660 31812 19669
rect 32036 19660 32088 19712
rect 33876 19660 33928 19712
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 1860 19363 1912 19372
rect 1860 19329 1869 19363
rect 1869 19329 1903 19363
rect 1903 19329 1912 19363
rect 1860 19320 1912 19329
rect 11796 19456 11848 19508
rect 12440 19456 12492 19508
rect 13360 19456 13412 19508
rect 15108 19456 15160 19508
rect 17316 19456 17368 19508
rect 18144 19499 18196 19508
rect 18144 19465 18153 19499
rect 18153 19465 18187 19499
rect 18187 19465 18196 19499
rect 26056 19499 26108 19508
rect 18144 19456 18196 19465
rect 12164 19388 12216 19440
rect 11980 19320 12032 19372
rect 12808 19388 12860 19440
rect 16120 19431 16172 19440
rect 16120 19397 16129 19431
rect 16129 19397 16163 19431
rect 16163 19397 16172 19431
rect 16120 19388 16172 19397
rect 12716 19363 12768 19372
rect 12716 19329 12725 19363
rect 12725 19329 12759 19363
rect 12759 19329 12768 19363
rect 13176 19363 13228 19372
rect 12716 19320 12768 19329
rect 13176 19329 13185 19363
rect 13185 19329 13219 19363
rect 13219 19329 13228 19363
rect 13176 19320 13228 19329
rect 13452 19363 13504 19372
rect 13452 19329 13486 19363
rect 13486 19329 13504 19363
rect 13452 19320 13504 19329
rect 15844 19320 15896 19372
rect 16580 19320 16632 19372
rect 16856 19320 16908 19372
rect 17592 19320 17644 19372
rect 2044 19295 2096 19304
rect 2044 19261 2053 19295
rect 2053 19261 2087 19295
rect 2087 19261 2096 19295
rect 2044 19252 2096 19261
rect 2780 19295 2832 19304
rect 2780 19261 2789 19295
rect 2789 19261 2823 19295
rect 2823 19261 2832 19295
rect 7932 19295 7984 19304
rect 2780 19252 2832 19261
rect 7932 19261 7941 19295
rect 7941 19261 7975 19295
rect 7975 19261 7984 19295
rect 7932 19252 7984 19261
rect 8208 19295 8260 19304
rect 8208 19261 8217 19295
rect 8217 19261 8251 19295
rect 8251 19261 8260 19295
rect 8208 19252 8260 19261
rect 19064 19388 19116 19440
rect 19432 19320 19484 19372
rect 20076 19388 20128 19440
rect 22652 19388 22704 19440
rect 22560 19320 22612 19372
rect 26056 19465 26065 19499
rect 26065 19465 26099 19499
rect 26099 19465 26108 19499
rect 26056 19456 26108 19465
rect 28632 19499 28684 19508
rect 28632 19465 28641 19499
rect 28641 19465 28675 19499
rect 28675 19465 28684 19499
rect 28632 19456 28684 19465
rect 30288 19499 30340 19508
rect 30288 19465 30297 19499
rect 30297 19465 30331 19499
rect 30331 19465 30340 19499
rect 30288 19456 30340 19465
rect 30656 19456 30708 19508
rect 31944 19456 31996 19508
rect 32404 19456 32456 19508
rect 33232 19456 33284 19508
rect 46756 19499 46808 19508
rect 46756 19465 46765 19499
rect 46765 19465 46799 19499
rect 46799 19465 46808 19499
rect 46756 19456 46808 19465
rect 23204 19431 23256 19440
rect 23204 19397 23213 19431
rect 23213 19397 23247 19431
rect 23247 19397 23256 19431
rect 23204 19388 23256 19397
rect 23940 19388 23992 19440
rect 21180 19252 21232 19304
rect 23940 19295 23992 19304
rect 23940 19261 23949 19295
rect 23949 19261 23983 19295
rect 23983 19261 23992 19295
rect 23940 19252 23992 19261
rect 24032 19252 24084 19304
rect 25412 19320 25464 19372
rect 28908 19363 28960 19372
rect 28908 19329 28917 19363
rect 28917 19329 28951 19363
rect 28951 19329 28960 19363
rect 28908 19320 28960 19329
rect 29092 19363 29144 19372
rect 29092 19329 29101 19363
rect 29101 19329 29135 19363
rect 29135 19329 29144 19363
rect 29092 19320 29144 19329
rect 29276 19363 29328 19372
rect 29276 19329 29285 19363
rect 29285 19329 29319 19363
rect 29319 19329 29328 19363
rect 29276 19320 29328 19329
rect 30012 19320 30064 19372
rect 31760 19388 31812 19440
rect 26424 19252 26476 19304
rect 31668 19320 31720 19372
rect 32312 19320 32364 19372
rect 47768 19295 47820 19304
rect 3516 19184 3568 19236
rect 12900 19184 12952 19236
rect 20720 19184 20772 19236
rect 12072 19159 12124 19168
rect 12072 19125 12081 19159
rect 12081 19125 12115 19159
rect 12115 19125 12124 19159
rect 12072 19116 12124 19125
rect 20536 19116 20588 19168
rect 22192 19116 22244 19168
rect 22284 19116 22336 19168
rect 28632 19184 28684 19236
rect 47768 19261 47777 19295
rect 47777 19261 47811 19295
rect 47811 19261 47820 19295
rect 47768 19252 47820 19261
rect 32220 19184 32272 19236
rect 24676 19116 24728 19168
rect 26608 19116 26660 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 2044 18912 2096 18964
rect 7932 18912 7984 18964
rect 9312 18912 9364 18964
rect 11796 18955 11848 18964
rect 9404 18844 9456 18896
rect 3792 18776 3844 18828
rect 7748 18776 7800 18828
rect 8300 18776 8352 18828
rect 7104 18751 7156 18760
rect 7104 18717 7113 18751
rect 7113 18717 7147 18751
rect 7147 18717 7156 18751
rect 7104 18708 7156 18717
rect 8024 18751 8076 18760
rect 8024 18717 8033 18751
rect 8033 18717 8067 18751
rect 8067 18717 8076 18751
rect 8024 18708 8076 18717
rect 8668 18708 8720 18760
rect 9588 18751 9640 18760
rect 9588 18717 9597 18751
rect 9597 18717 9631 18751
rect 9631 18717 9640 18751
rect 9588 18708 9640 18717
rect 11796 18921 11805 18955
rect 11805 18921 11839 18955
rect 11839 18921 11848 18955
rect 11796 18912 11848 18921
rect 11980 18912 12032 18964
rect 13360 18912 13412 18964
rect 17500 18912 17552 18964
rect 25412 18912 25464 18964
rect 26424 18955 26476 18964
rect 26424 18921 26433 18955
rect 26433 18921 26467 18955
rect 26467 18921 26476 18955
rect 26424 18912 26476 18921
rect 29092 18912 29144 18964
rect 30196 18912 30248 18964
rect 32312 18912 32364 18964
rect 15660 18844 15712 18896
rect 25872 18844 25924 18896
rect 26240 18844 26292 18896
rect 12256 18819 12308 18828
rect 12256 18785 12265 18819
rect 12265 18785 12299 18819
rect 12299 18785 12308 18819
rect 12256 18776 12308 18785
rect 10416 18751 10468 18760
rect 10416 18717 10425 18751
rect 10425 18717 10459 18751
rect 10459 18717 10468 18751
rect 10416 18708 10468 18717
rect 12072 18708 12124 18760
rect 12440 18708 12492 18760
rect 15752 18751 15804 18760
rect 15752 18717 15761 18751
rect 15761 18717 15795 18751
rect 15795 18717 15804 18751
rect 15752 18708 15804 18717
rect 18052 18776 18104 18828
rect 22652 18776 22704 18828
rect 6828 18572 6880 18624
rect 8944 18615 8996 18624
rect 8944 18581 8953 18615
rect 8953 18581 8987 18615
rect 8987 18581 8996 18615
rect 8944 18572 8996 18581
rect 10600 18640 10652 18692
rect 18144 18708 18196 18760
rect 22468 18751 22520 18760
rect 22468 18717 22477 18751
rect 22477 18717 22511 18751
rect 22511 18717 22520 18751
rect 22468 18708 22520 18717
rect 24676 18708 24728 18760
rect 24952 18708 25004 18760
rect 25412 18708 25464 18760
rect 26148 18751 26200 18760
rect 25136 18683 25188 18692
rect 25136 18649 25145 18683
rect 25145 18649 25179 18683
rect 25179 18649 25188 18683
rect 25136 18640 25188 18649
rect 25780 18640 25832 18692
rect 26148 18717 26157 18751
rect 26157 18717 26191 18751
rect 26191 18717 26200 18751
rect 26148 18708 26200 18717
rect 28908 18844 28960 18896
rect 28724 18776 28776 18828
rect 47308 18819 47360 18828
rect 27804 18708 27856 18760
rect 31852 18751 31904 18760
rect 31852 18717 31861 18751
rect 31861 18717 31895 18751
rect 31895 18717 31904 18751
rect 31852 18708 31904 18717
rect 11888 18572 11940 18624
rect 23664 18572 23716 18624
rect 24400 18572 24452 18624
rect 24584 18572 24636 18624
rect 26608 18640 26660 18692
rect 27988 18683 28040 18692
rect 27988 18649 27997 18683
rect 27997 18649 28031 18683
rect 28031 18649 28040 18683
rect 27988 18640 28040 18649
rect 28632 18683 28684 18692
rect 28632 18649 28641 18683
rect 28641 18649 28675 18683
rect 28675 18649 28684 18683
rect 28632 18640 28684 18649
rect 29920 18640 29972 18692
rect 32036 18751 32088 18760
rect 32036 18717 32045 18751
rect 32045 18717 32079 18751
rect 32079 18717 32088 18751
rect 32036 18708 32088 18717
rect 32220 18751 32272 18760
rect 32220 18717 32229 18751
rect 32229 18717 32263 18751
rect 32263 18717 32272 18751
rect 32220 18708 32272 18717
rect 32588 18708 32640 18760
rect 47308 18785 47317 18819
rect 47317 18785 47351 18819
rect 47351 18785 47360 18819
rect 47308 18776 47360 18785
rect 46204 18708 46256 18760
rect 29276 18572 29328 18624
rect 31944 18572 31996 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 7840 18368 7892 18420
rect 6828 18343 6880 18352
rect 6828 18309 6837 18343
rect 6837 18309 6871 18343
rect 6871 18309 6880 18343
rect 6828 18300 6880 18309
rect 2688 18275 2740 18284
rect 2688 18241 2697 18275
rect 2697 18241 2731 18275
rect 2731 18241 2740 18275
rect 2688 18232 2740 18241
rect 22100 18368 22152 18420
rect 24676 18368 24728 18420
rect 8944 18300 8996 18352
rect 10600 18343 10652 18352
rect 10600 18309 10609 18343
rect 10609 18309 10643 18343
rect 10643 18309 10652 18343
rect 10600 18300 10652 18309
rect 10968 18343 11020 18352
rect 10968 18309 10977 18343
rect 10977 18309 11011 18343
rect 11011 18309 11020 18343
rect 10968 18300 11020 18309
rect 2320 18164 2372 18216
rect 10876 18232 10928 18284
rect 11980 18232 12032 18284
rect 7840 18207 7892 18216
rect 7840 18173 7849 18207
rect 7849 18173 7883 18207
rect 7883 18173 7892 18207
rect 7840 18164 7892 18173
rect 11796 18164 11848 18216
rect 12256 18278 12308 18284
rect 12256 18244 12265 18278
rect 12265 18244 12299 18278
rect 12299 18244 12308 18278
rect 12440 18275 12492 18284
rect 12256 18232 12308 18244
rect 12440 18241 12449 18275
rect 12449 18241 12483 18275
rect 12483 18241 12492 18275
rect 12440 18232 12492 18241
rect 12900 18232 12952 18284
rect 15108 18300 15160 18352
rect 15660 18343 15712 18352
rect 15660 18309 15669 18343
rect 15669 18309 15703 18343
rect 15703 18309 15712 18343
rect 15660 18300 15712 18309
rect 17592 18300 17644 18352
rect 19432 18300 19484 18352
rect 25780 18368 25832 18420
rect 3148 18096 3200 18148
rect 9588 18096 9640 18148
rect 14188 18232 14240 18284
rect 14556 18232 14608 18284
rect 15844 18232 15896 18284
rect 17960 18232 18012 18284
rect 13268 18096 13320 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2136 18071 2188 18080
rect 2136 18037 2145 18071
rect 2145 18037 2179 18071
rect 2179 18037 2188 18071
rect 2136 18028 2188 18037
rect 2872 18028 2924 18080
rect 8760 18028 8812 18080
rect 11796 18071 11848 18080
rect 11796 18037 11805 18071
rect 11805 18037 11839 18071
rect 11839 18037 11848 18071
rect 11796 18028 11848 18037
rect 11888 18028 11940 18080
rect 12900 18028 12952 18080
rect 13452 18071 13504 18080
rect 13452 18037 13461 18071
rect 13461 18037 13495 18071
rect 13495 18037 13504 18071
rect 13452 18028 13504 18037
rect 13912 18096 13964 18148
rect 14004 18096 14056 18148
rect 18420 18096 18472 18148
rect 18788 18232 18840 18284
rect 20628 18232 20680 18284
rect 21180 18232 21232 18284
rect 23204 18232 23256 18284
rect 23480 18232 23532 18284
rect 25872 18300 25924 18352
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 25320 18232 25372 18284
rect 26240 18232 26292 18284
rect 27620 18275 27672 18284
rect 27620 18241 27629 18275
rect 27629 18241 27663 18275
rect 27663 18241 27672 18275
rect 27620 18232 27672 18241
rect 28264 18232 28316 18284
rect 24032 18164 24084 18216
rect 19340 18096 19392 18148
rect 22928 18096 22980 18148
rect 24676 18096 24728 18148
rect 15384 18028 15436 18080
rect 18144 18028 18196 18080
rect 18604 18028 18656 18080
rect 23296 18028 23348 18080
rect 23848 18071 23900 18080
rect 23848 18037 23857 18071
rect 23857 18037 23891 18071
rect 23891 18037 23900 18071
rect 23848 18028 23900 18037
rect 24032 18071 24084 18080
rect 24032 18037 24041 18071
rect 24041 18037 24075 18071
rect 24075 18037 24084 18071
rect 24032 18028 24084 18037
rect 26056 18164 26108 18216
rect 25320 18028 25372 18080
rect 29000 18071 29052 18080
rect 29000 18037 29009 18071
rect 29009 18037 29043 18071
rect 29043 18037 29052 18071
rect 29000 18028 29052 18037
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 8300 17824 8352 17876
rect 9312 17756 9364 17808
rect 1584 17688 1636 17740
rect 2780 17731 2832 17740
rect 2780 17697 2789 17731
rect 2789 17697 2823 17731
rect 2823 17697 2832 17731
rect 2780 17688 2832 17697
rect 7932 17620 7984 17672
rect 2136 17552 2188 17604
rect 7380 17595 7432 17604
rect 7380 17561 7389 17595
rect 7389 17561 7423 17595
rect 7423 17561 7432 17595
rect 7380 17552 7432 17561
rect 10876 17824 10928 17876
rect 14004 17824 14056 17876
rect 20628 17867 20680 17876
rect 9588 17663 9640 17672
rect 9588 17629 9597 17663
rect 9597 17629 9631 17663
rect 9631 17629 9640 17663
rect 9588 17620 9640 17629
rect 10416 17620 10468 17672
rect 8760 17484 8812 17536
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 9496 17552 9548 17604
rect 11796 17620 11848 17672
rect 13176 17756 13228 17808
rect 13912 17756 13964 17808
rect 17592 17799 17644 17808
rect 17592 17765 17601 17799
rect 17601 17765 17635 17799
rect 17635 17765 17644 17799
rect 17592 17756 17644 17765
rect 9220 17484 9272 17536
rect 12992 17620 13044 17672
rect 13268 17620 13320 17672
rect 15752 17620 15804 17672
rect 18512 17756 18564 17808
rect 14372 17595 14424 17604
rect 14372 17561 14381 17595
rect 14381 17561 14415 17595
rect 14415 17561 14424 17595
rect 14372 17552 14424 17561
rect 17684 17552 17736 17604
rect 15476 17484 15528 17536
rect 16764 17484 16816 17536
rect 18236 17620 18288 17672
rect 20628 17833 20637 17867
rect 20637 17833 20671 17867
rect 20671 17833 20680 17867
rect 20628 17824 20680 17833
rect 19248 17731 19300 17740
rect 19248 17697 19257 17731
rect 19257 17697 19291 17731
rect 19291 17697 19300 17731
rect 19248 17688 19300 17697
rect 18604 17552 18656 17604
rect 18788 17552 18840 17604
rect 18420 17484 18472 17536
rect 18512 17484 18564 17536
rect 20812 17620 20864 17672
rect 22468 17824 22520 17876
rect 23020 17824 23072 17876
rect 24124 17824 24176 17876
rect 22652 17756 22704 17808
rect 23480 17756 23532 17808
rect 22928 17688 22980 17740
rect 23388 17688 23440 17740
rect 26148 17824 26200 17876
rect 26884 17824 26936 17876
rect 24952 17756 25004 17808
rect 28080 17756 28132 17808
rect 22100 17663 22152 17672
rect 22100 17629 22109 17663
rect 22109 17629 22143 17663
rect 22143 17629 22152 17663
rect 22100 17620 22152 17629
rect 22468 17620 22520 17672
rect 20628 17552 20680 17604
rect 22652 17552 22704 17604
rect 23296 17620 23348 17672
rect 24584 17552 24636 17604
rect 20076 17484 20128 17536
rect 20352 17484 20404 17536
rect 22284 17484 22336 17536
rect 22468 17484 22520 17536
rect 22928 17527 22980 17536
rect 22928 17493 22937 17527
rect 22937 17493 22971 17527
rect 22971 17493 22980 17527
rect 22928 17484 22980 17493
rect 23020 17484 23072 17536
rect 25136 17620 25188 17672
rect 25872 17663 25924 17672
rect 25872 17629 25881 17663
rect 25881 17629 25915 17663
rect 25915 17629 25924 17663
rect 25872 17620 25924 17629
rect 25320 17552 25372 17604
rect 27436 17620 27488 17672
rect 27620 17663 27672 17672
rect 27620 17629 27629 17663
rect 27629 17629 27663 17663
rect 27663 17629 27672 17663
rect 27620 17620 27672 17629
rect 24952 17527 25004 17536
rect 24952 17493 24961 17527
rect 24961 17493 24995 17527
rect 24995 17493 25004 17527
rect 24952 17484 25004 17493
rect 27896 17688 27948 17740
rect 29184 17688 29236 17740
rect 30012 17731 30064 17740
rect 30012 17697 30021 17731
rect 30021 17697 30055 17731
rect 30055 17697 30064 17731
rect 30012 17688 30064 17697
rect 28172 17620 28224 17672
rect 28448 17663 28500 17672
rect 28448 17629 28457 17663
rect 28457 17629 28491 17663
rect 28491 17629 28500 17663
rect 28448 17620 28500 17629
rect 29276 17620 29328 17672
rect 46296 17620 46348 17672
rect 29000 17552 29052 17604
rect 28356 17484 28408 17536
rect 28724 17527 28776 17536
rect 28724 17493 28733 17527
rect 28733 17493 28767 17527
rect 28767 17493 28776 17527
rect 28724 17484 28776 17493
rect 29828 17484 29880 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 7932 17280 7984 17332
rect 9312 17280 9364 17332
rect 2872 17212 2924 17264
rect 7380 17212 7432 17264
rect 7840 17187 7892 17196
rect 7840 17153 7849 17187
rect 7849 17153 7883 17187
rect 7883 17153 7892 17187
rect 7840 17144 7892 17153
rect 8944 17144 8996 17196
rect 13452 17187 13504 17196
rect 13452 17153 13486 17187
rect 13486 17153 13504 17187
rect 13452 17144 13504 17153
rect 15568 17212 15620 17264
rect 1400 17119 1452 17128
rect 1400 17085 1409 17119
rect 1409 17085 1443 17119
rect 1443 17085 1452 17119
rect 1400 17076 1452 17085
rect 2780 17119 2832 17128
rect 2780 17085 2789 17119
rect 2789 17085 2823 17119
rect 2823 17085 2832 17119
rect 3884 17119 3936 17128
rect 2780 17076 2832 17085
rect 3884 17085 3893 17119
rect 3893 17085 3927 17119
rect 3927 17085 3936 17119
rect 3884 17076 3936 17085
rect 4068 17076 4120 17128
rect 13176 17119 13228 17128
rect 13176 17085 13185 17119
rect 13185 17085 13219 17119
rect 13219 17085 13228 17119
rect 13176 17076 13228 17085
rect 15016 17119 15068 17128
rect 15016 17085 15025 17119
rect 15025 17085 15059 17119
rect 15059 17085 15068 17119
rect 15016 17076 15068 17085
rect 15476 17187 15528 17196
rect 15476 17153 15485 17187
rect 15485 17153 15519 17187
rect 15519 17153 15528 17187
rect 15476 17144 15528 17153
rect 15660 17187 15712 17196
rect 15660 17153 15669 17187
rect 15669 17153 15703 17187
rect 15703 17153 15712 17187
rect 16764 17187 16816 17196
rect 15660 17144 15712 17153
rect 16764 17153 16773 17187
rect 16773 17153 16807 17187
rect 16807 17153 16816 17187
rect 16764 17144 16816 17153
rect 16948 17187 17000 17196
rect 16948 17153 16957 17187
rect 16957 17153 16991 17187
rect 16991 17153 17000 17187
rect 16948 17144 17000 17153
rect 17408 17187 17460 17196
rect 17408 17153 17417 17187
rect 17417 17153 17451 17187
rect 17451 17153 17460 17187
rect 17408 17144 17460 17153
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 18420 17212 18472 17264
rect 18604 17280 18656 17332
rect 19248 17280 19300 17332
rect 24860 17280 24912 17332
rect 26332 17323 26384 17332
rect 26332 17289 26341 17323
rect 26341 17289 26375 17323
rect 26375 17289 26384 17323
rect 26332 17280 26384 17289
rect 30012 17323 30064 17332
rect 30012 17289 30021 17323
rect 30021 17289 30055 17323
rect 30055 17289 30064 17323
rect 30012 17280 30064 17289
rect 18144 17144 18196 17196
rect 19616 17144 19668 17196
rect 16580 17076 16632 17128
rect 14556 17051 14608 17060
rect 14556 17017 14565 17051
rect 14565 17017 14599 17051
rect 14599 17017 14608 17051
rect 14556 17008 14608 17017
rect 14832 17008 14884 17060
rect 1768 16940 1820 16992
rect 9312 16940 9364 16992
rect 15108 17008 15160 17060
rect 15660 17008 15712 17060
rect 19432 17051 19484 17060
rect 19432 17017 19441 17051
rect 19441 17017 19475 17051
rect 19475 17017 19484 17051
rect 22468 17144 22520 17196
rect 22652 17076 22704 17128
rect 23296 17212 23348 17264
rect 23388 17212 23440 17264
rect 27620 17212 27672 17264
rect 28724 17212 28776 17264
rect 29460 17212 29512 17264
rect 31024 17212 31076 17264
rect 46388 17212 46440 17264
rect 23204 17187 23256 17196
rect 23204 17153 23213 17187
rect 23213 17153 23247 17187
rect 23247 17153 23256 17187
rect 23664 17187 23716 17196
rect 23204 17144 23256 17153
rect 23664 17153 23673 17187
rect 23673 17153 23707 17187
rect 23707 17153 23716 17187
rect 23664 17144 23716 17153
rect 24032 17144 24084 17196
rect 19432 17008 19484 17017
rect 22468 17008 22520 17060
rect 18420 16940 18472 16992
rect 18788 16940 18840 16992
rect 20628 16940 20680 16992
rect 22376 16940 22428 16992
rect 23388 17076 23440 17128
rect 23296 17008 23348 17060
rect 23664 17008 23716 17060
rect 26056 17144 26108 17196
rect 28172 17144 28224 17196
rect 28908 17187 28960 17196
rect 28908 17153 28917 17187
rect 28917 17153 28951 17187
rect 28951 17153 28960 17187
rect 28908 17144 28960 17153
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 31668 17144 31720 17196
rect 33508 17144 33560 17196
rect 47216 17144 47268 17196
rect 24584 17076 24636 17128
rect 24216 17008 24268 17060
rect 25872 17076 25924 17128
rect 27436 17119 27488 17128
rect 27436 17085 27445 17119
rect 27445 17085 27479 17119
rect 27479 17085 27488 17119
rect 27436 17076 27488 17085
rect 28448 17076 28500 17128
rect 30104 17119 30156 17128
rect 30104 17085 30113 17119
rect 30113 17085 30147 17119
rect 30147 17085 30156 17119
rect 30104 17076 30156 17085
rect 30288 17119 30340 17128
rect 30288 17085 30297 17119
rect 30297 17085 30331 17119
rect 30331 17085 30340 17119
rect 30288 17076 30340 17085
rect 30012 17008 30064 17060
rect 29184 16940 29236 16992
rect 29736 16940 29788 16992
rect 32128 16940 32180 16992
rect 33048 16940 33100 16992
rect 47032 16983 47084 16992
rect 47032 16949 47041 16983
rect 47041 16949 47075 16983
rect 47075 16949 47084 16983
rect 47032 16940 47084 16949
rect 47676 16983 47728 16992
rect 47676 16949 47685 16983
rect 47685 16949 47719 16983
rect 47719 16949 47728 16983
rect 47676 16940 47728 16949
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 1400 16736 1452 16788
rect 3884 16779 3936 16788
rect 3884 16745 3893 16779
rect 3893 16745 3927 16779
rect 3927 16745 3936 16779
rect 3884 16736 3936 16745
rect 13176 16668 13228 16720
rect 13728 16668 13780 16720
rect 16948 16736 17000 16788
rect 17500 16736 17552 16788
rect 17592 16736 17644 16788
rect 18788 16668 18840 16720
rect 19340 16736 19392 16788
rect 22652 16736 22704 16788
rect 20076 16668 20128 16720
rect 22100 16668 22152 16720
rect 1860 16575 1912 16584
rect 1860 16541 1869 16575
rect 1869 16541 1903 16575
rect 1903 16541 1912 16575
rect 1860 16532 1912 16541
rect 8024 16600 8076 16652
rect 10876 16600 10928 16652
rect 11428 16643 11480 16652
rect 11428 16609 11437 16643
rect 11437 16609 11471 16643
rect 11471 16609 11480 16643
rect 11428 16600 11480 16609
rect 13912 16600 13964 16652
rect 15384 16643 15436 16652
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 15384 16609 15393 16643
rect 15393 16609 15427 16643
rect 15427 16609 15436 16643
rect 15384 16600 15436 16609
rect 19340 16600 19392 16652
rect 19616 16600 19668 16652
rect 22284 16600 22336 16652
rect 15108 16532 15160 16584
rect 11612 16464 11664 16516
rect 14832 16464 14884 16516
rect 20 16396 72 16448
rect 11428 16396 11480 16448
rect 16580 16396 16632 16448
rect 17592 16532 17644 16584
rect 20260 16532 20312 16584
rect 20628 16575 20680 16584
rect 20628 16541 20637 16575
rect 20637 16541 20671 16575
rect 20671 16541 20680 16575
rect 20628 16532 20680 16541
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 17684 16464 17736 16516
rect 18696 16507 18748 16516
rect 18696 16473 18705 16507
rect 18705 16473 18739 16507
rect 18739 16473 18748 16507
rect 18696 16464 18748 16473
rect 19432 16507 19484 16516
rect 19432 16473 19441 16507
rect 19441 16473 19475 16507
rect 19475 16473 19484 16507
rect 19432 16464 19484 16473
rect 19524 16464 19576 16516
rect 22192 16439 22244 16448
rect 22192 16405 22201 16439
rect 22201 16405 22235 16439
rect 22235 16405 22244 16439
rect 22192 16396 22244 16405
rect 22468 16600 22520 16652
rect 23020 16668 23072 16720
rect 23848 16736 23900 16788
rect 25136 16736 25188 16788
rect 25964 16736 26016 16788
rect 28264 16779 28316 16788
rect 28264 16745 28273 16779
rect 28273 16745 28307 16779
rect 28307 16745 28316 16779
rect 28264 16736 28316 16745
rect 24860 16668 24912 16720
rect 22928 16600 22980 16652
rect 23480 16643 23532 16652
rect 23480 16609 23489 16643
rect 23489 16609 23523 16643
rect 23523 16609 23532 16643
rect 23480 16600 23532 16609
rect 26424 16600 26476 16652
rect 27160 16600 27212 16652
rect 29736 16668 29788 16720
rect 30748 16668 30800 16720
rect 25320 16532 25372 16584
rect 22560 16507 22612 16516
rect 22560 16473 22569 16507
rect 22569 16473 22603 16507
rect 22603 16473 22612 16507
rect 22560 16464 22612 16473
rect 23296 16464 23348 16516
rect 23480 16464 23532 16516
rect 24492 16464 24544 16516
rect 26056 16464 26108 16516
rect 26976 16532 27028 16584
rect 27252 16532 27304 16584
rect 27620 16532 27672 16584
rect 29092 16600 29144 16652
rect 31668 16736 31720 16788
rect 33508 16779 33560 16788
rect 33508 16745 33517 16779
rect 33517 16745 33551 16779
rect 33551 16745 33560 16779
rect 33508 16736 33560 16745
rect 32128 16668 32180 16720
rect 22652 16396 22704 16448
rect 23020 16396 23072 16448
rect 24400 16396 24452 16448
rect 25688 16396 25740 16448
rect 26424 16396 26476 16448
rect 28356 16532 28408 16584
rect 28724 16464 28776 16516
rect 29828 16575 29880 16584
rect 29828 16541 29837 16575
rect 29837 16541 29871 16575
rect 29871 16541 29880 16575
rect 29828 16532 29880 16541
rect 30012 16575 30064 16584
rect 30012 16541 30021 16575
rect 30021 16541 30055 16575
rect 30055 16541 30064 16575
rect 30012 16532 30064 16541
rect 33048 16643 33100 16652
rect 33048 16609 33057 16643
rect 33057 16609 33091 16643
rect 33091 16609 33100 16643
rect 33048 16600 33100 16609
rect 46296 16643 46348 16652
rect 46296 16609 46305 16643
rect 46305 16609 46339 16643
rect 46339 16609 46348 16643
rect 46296 16600 46348 16609
rect 48136 16643 48188 16652
rect 48136 16609 48145 16643
rect 48145 16609 48179 16643
rect 48179 16609 48188 16643
rect 48136 16600 48188 16609
rect 29736 16464 29788 16516
rect 30104 16507 30156 16516
rect 30104 16473 30113 16507
rect 30113 16473 30147 16507
rect 30147 16473 30156 16507
rect 30104 16464 30156 16473
rect 30748 16464 30800 16516
rect 30932 16396 30984 16448
rect 31576 16532 31628 16584
rect 32956 16575 33008 16584
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 32956 16532 33008 16541
rect 31392 16464 31444 16516
rect 47676 16464 47728 16516
rect 32312 16439 32364 16448
rect 32312 16405 32321 16439
rect 32321 16405 32355 16439
rect 32355 16405 32364 16439
rect 32312 16396 32364 16405
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 11612 16235 11664 16244
rect 11612 16201 11621 16235
rect 11621 16201 11655 16235
rect 11655 16201 11664 16235
rect 11612 16192 11664 16201
rect 17500 16235 17552 16244
rect 17500 16201 17509 16235
rect 17509 16201 17543 16235
rect 17543 16201 17552 16235
rect 17500 16192 17552 16201
rect 18420 16192 18472 16244
rect 22100 16192 22152 16244
rect 24400 16192 24452 16244
rect 29000 16235 29052 16244
rect 24032 16167 24084 16176
rect 11520 16099 11572 16108
rect 11520 16065 11529 16099
rect 11529 16065 11563 16099
rect 11563 16065 11572 16099
rect 24032 16133 24041 16167
rect 24041 16133 24075 16167
rect 24075 16133 24084 16167
rect 24032 16124 24084 16133
rect 24676 16124 24728 16176
rect 24952 16124 25004 16176
rect 29000 16201 29009 16235
rect 29009 16201 29043 16235
rect 29043 16201 29052 16235
rect 29000 16192 29052 16201
rect 28448 16124 28500 16176
rect 29184 16124 29236 16176
rect 13728 16099 13780 16108
rect 11520 16056 11572 16065
rect 13728 16065 13737 16099
rect 13737 16065 13771 16099
rect 13771 16065 13780 16099
rect 13728 16056 13780 16065
rect 15016 16056 15068 16108
rect 17316 16099 17368 16108
rect 17316 16065 17325 16099
rect 17325 16065 17359 16099
rect 17359 16065 17368 16099
rect 17316 16056 17368 16065
rect 17408 16056 17460 16108
rect 17868 15988 17920 16040
rect 18788 16099 18840 16108
rect 18788 16065 18797 16099
rect 18797 16065 18831 16099
rect 18831 16065 18840 16099
rect 18788 16056 18840 16065
rect 19248 16099 19300 16108
rect 19248 16065 19257 16099
rect 19257 16065 19291 16099
rect 19291 16065 19300 16099
rect 19248 16056 19300 16065
rect 22192 16056 22244 16108
rect 22652 16099 22704 16108
rect 22652 16065 22661 16099
rect 22661 16065 22695 16099
rect 22695 16065 22704 16099
rect 22652 16056 22704 16065
rect 23020 16056 23072 16108
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 20628 15963 20680 15972
rect 20628 15929 20637 15963
rect 20637 15929 20671 15963
rect 20671 15929 20680 15963
rect 22928 16031 22980 16040
rect 22928 15997 22937 16031
rect 22937 15997 22971 16031
rect 22971 15997 22980 16031
rect 22928 15988 22980 15997
rect 20628 15920 20680 15929
rect 15108 15895 15160 15904
rect 15108 15861 15117 15895
rect 15117 15861 15151 15895
rect 15151 15861 15160 15895
rect 15108 15852 15160 15861
rect 17132 15895 17184 15904
rect 17132 15861 17141 15895
rect 17141 15861 17175 15895
rect 17175 15861 17184 15895
rect 17132 15852 17184 15861
rect 22284 15852 22336 15904
rect 24124 15920 24176 15972
rect 25044 16056 25096 16108
rect 26976 16099 27028 16108
rect 26976 16065 26985 16099
rect 26985 16065 27019 16099
rect 27019 16065 27028 16099
rect 26976 16056 27028 16065
rect 27160 16099 27212 16108
rect 27160 16065 27169 16099
rect 27169 16065 27203 16099
rect 27203 16065 27212 16099
rect 27160 16056 27212 16065
rect 27804 16099 27856 16108
rect 27804 16065 27813 16099
rect 27813 16065 27847 16099
rect 27847 16065 27856 16099
rect 27804 16056 27856 16065
rect 28080 16099 28132 16108
rect 28080 16065 28089 16099
rect 28089 16065 28123 16099
rect 28123 16065 28132 16099
rect 28080 16056 28132 16065
rect 30196 16192 30248 16244
rect 30564 16192 30616 16244
rect 30840 16167 30892 16176
rect 30840 16133 30849 16167
rect 30849 16133 30883 16167
rect 30883 16133 30892 16167
rect 30840 16124 30892 16133
rect 33048 16124 33100 16176
rect 29460 16099 29512 16108
rect 29460 16065 29469 16099
rect 29469 16065 29503 16099
rect 29503 16065 29512 16099
rect 29460 16056 29512 16065
rect 31392 16056 31444 16108
rect 32312 16099 32364 16108
rect 32312 16065 32321 16099
rect 32321 16065 32355 16099
rect 32355 16065 32364 16099
rect 32312 16056 32364 16065
rect 32404 16099 32456 16108
rect 32404 16065 32413 16099
rect 32413 16065 32447 16099
rect 32447 16065 32456 16099
rect 32404 16056 32456 16065
rect 47216 16056 47268 16108
rect 24860 15988 24912 16040
rect 25320 15988 25372 16040
rect 29552 15988 29604 16040
rect 31024 16031 31076 16040
rect 25504 15920 25556 15972
rect 27896 15920 27948 15972
rect 31024 15997 31033 16031
rect 31033 15997 31067 16031
rect 31067 15997 31076 16031
rect 31024 15988 31076 15997
rect 25596 15895 25648 15904
rect 25596 15861 25605 15895
rect 25605 15861 25639 15895
rect 25639 15861 25648 15895
rect 25596 15852 25648 15861
rect 26332 15852 26384 15904
rect 29184 15852 29236 15904
rect 30380 15852 30432 15904
rect 31576 15852 31628 15904
rect 32128 15895 32180 15904
rect 32128 15861 32137 15895
rect 32137 15861 32171 15895
rect 32171 15861 32180 15895
rect 32128 15852 32180 15861
rect 32312 15852 32364 15904
rect 46480 15852 46532 15904
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 17408 15648 17460 15700
rect 22468 15691 22520 15700
rect 22468 15657 22477 15691
rect 22477 15657 22511 15691
rect 22511 15657 22520 15691
rect 22468 15648 22520 15657
rect 22928 15691 22980 15700
rect 22928 15657 22937 15691
rect 22937 15657 22971 15691
rect 22971 15657 22980 15691
rect 22928 15648 22980 15657
rect 24768 15648 24820 15700
rect 25596 15648 25648 15700
rect 26976 15648 27028 15700
rect 28908 15648 28960 15700
rect 14372 15580 14424 15632
rect 15108 15580 15160 15632
rect 17868 15580 17920 15632
rect 12348 15555 12400 15564
rect 12348 15521 12357 15555
rect 12357 15521 12391 15555
rect 12391 15521 12400 15555
rect 12348 15512 12400 15521
rect 19248 15512 19300 15564
rect 12900 15487 12952 15496
rect 12900 15453 12909 15487
rect 12909 15453 12943 15487
rect 12943 15453 12952 15487
rect 12900 15444 12952 15453
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 28172 15580 28224 15632
rect 30012 15580 30064 15632
rect 25320 15555 25372 15564
rect 25320 15521 25329 15555
rect 25329 15521 25363 15555
rect 25363 15521 25372 15555
rect 25320 15512 25372 15521
rect 26056 15512 26108 15564
rect 30288 15648 30340 15700
rect 30932 15580 30984 15632
rect 31852 15580 31904 15632
rect 23112 15487 23164 15496
rect 10784 15419 10836 15428
rect 10784 15385 10793 15419
rect 10793 15385 10827 15419
rect 10827 15385 10836 15419
rect 10784 15376 10836 15385
rect 17132 15376 17184 15428
rect 18788 15376 18840 15428
rect 23112 15453 23121 15487
rect 23121 15453 23155 15487
rect 23155 15453 23164 15487
rect 23112 15444 23164 15453
rect 23296 15487 23348 15496
rect 23296 15453 23305 15487
rect 23305 15453 23339 15487
rect 23339 15453 23348 15487
rect 23296 15444 23348 15453
rect 24492 15487 24544 15496
rect 22100 15376 22152 15428
rect 12624 15308 12676 15360
rect 20996 15308 21048 15360
rect 24492 15453 24501 15487
rect 24501 15453 24535 15487
rect 24535 15453 24544 15487
rect 24492 15444 24544 15453
rect 24952 15444 25004 15496
rect 25504 15487 25556 15496
rect 25504 15453 25513 15487
rect 25513 15453 25547 15487
rect 25547 15453 25556 15487
rect 25504 15444 25556 15453
rect 27160 15444 27212 15496
rect 24124 15376 24176 15428
rect 26332 15419 26384 15428
rect 26332 15385 26357 15419
rect 26357 15385 26384 15419
rect 27896 15419 27948 15428
rect 26332 15376 26384 15385
rect 27896 15385 27905 15419
rect 27905 15385 27939 15419
rect 27939 15385 27948 15419
rect 27896 15376 27948 15385
rect 28448 15444 28500 15496
rect 28724 15487 28776 15496
rect 28724 15453 28733 15487
rect 28733 15453 28767 15487
rect 28767 15453 28776 15487
rect 28724 15444 28776 15453
rect 30012 15444 30064 15496
rect 30196 15487 30248 15496
rect 30196 15453 30205 15487
rect 30205 15453 30239 15487
rect 30239 15453 30248 15487
rect 30196 15444 30248 15453
rect 30748 15512 30800 15564
rect 32956 15580 33008 15632
rect 47032 15580 47084 15632
rect 46480 15555 46532 15564
rect 46480 15521 46489 15555
rect 46489 15521 46523 15555
rect 46523 15521 46532 15555
rect 46480 15512 46532 15521
rect 48136 15555 48188 15564
rect 48136 15521 48145 15555
rect 48145 15521 48179 15555
rect 48179 15521 48188 15555
rect 48136 15512 48188 15521
rect 30840 15487 30892 15496
rect 30840 15453 30849 15487
rect 30849 15453 30883 15487
rect 30883 15453 30892 15487
rect 30840 15444 30892 15453
rect 29644 15376 29696 15428
rect 31760 15487 31812 15496
rect 31760 15453 31769 15487
rect 31769 15453 31803 15487
rect 31803 15453 31812 15487
rect 31760 15444 31812 15453
rect 31944 15487 31996 15496
rect 31944 15453 31953 15487
rect 31953 15453 31987 15487
rect 31987 15453 31996 15487
rect 31944 15444 31996 15453
rect 32404 15444 32456 15496
rect 33324 15444 33376 15496
rect 33968 15444 34020 15496
rect 26056 15308 26108 15360
rect 26516 15351 26568 15360
rect 26516 15317 26525 15351
rect 26525 15317 26559 15351
rect 26559 15317 26568 15351
rect 26516 15308 26568 15317
rect 26884 15308 26936 15360
rect 29460 15308 29512 15360
rect 30472 15308 30524 15360
rect 32496 15351 32548 15360
rect 32496 15317 32505 15351
rect 32505 15317 32539 15351
rect 32539 15317 32548 15351
rect 32496 15308 32548 15317
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 10784 15147 10836 15156
rect 10784 15113 10793 15147
rect 10793 15113 10827 15147
rect 10827 15113 10836 15147
rect 10784 15104 10836 15113
rect 22100 15147 22152 15156
rect 22100 15113 22109 15147
rect 22109 15113 22143 15147
rect 22143 15113 22152 15147
rect 22100 15104 22152 15113
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 23112 15036 23164 15088
rect 22284 15011 22336 15020
rect 22284 14977 22293 15011
rect 22293 14977 22327 15011
rect 22327 14977 22336 15011
rect 22284 14968 22336 14977
rect 22468 14968 22520 15020
rect 24032 15011 24084 15020
rect 24032 14977 24041 15011
rect 24041 14977 24075 15011
rect 24075 14977 24084 15011
rect 24032 14968 24084 14977
rect 25504 15104 25556 15156
rect 27896 15104 27948 15156
rect 27436 15036 27488 15088
rect 30380 15104 30432 15156
rect 31760 15104 31812 15156
rect 33968 15147 34020 15156
rect 33968 15113 33977 15147
rect 33977 15113 34011 15147
rect 34011 15113 34020 15147
rect 33968 15104 34020 15113
rect 47860 15104 47912 15156
rect 29000 15036 29052 15088
rect 24400 14968 24452 15020
rect 24584 14968 24636 15020
rect 24860 14968 24912 15020
rect 26148 14968 26200 15020
rect 26516 14968 26568 15020
rect 27528 14968 27580 15020
rect 29644 15011 29696 15020
rect 29644 14977 29653 15011
rect 29653 14977 29687 15011
rect 29687 14977 29696 15011
rect 29644 14968 29696 14977
rect 19432 14900 19484 14952
rect 20996 14900 21048 14952
rect 26240 14900 26292 14952
rect 29552 14943 29604 14952
rect 29552 14909 29561 14943
rect 29561 14909 29595 14943
rect 29595 14909 29604 14943
rect 29552 14900 29604 14909
rect 32496 15036 32548 15088
rect 30472 15011 30524 15020
rect 30472 14977 30481 15011
rect 30481 14977 30515 15011
rect 30515 14977 30524 15011
rect 30472 14968 30524 14977
rect 30564 15011 30616 15020
rect 30564 14977 30573 15011
rect 30573 14977 30607 15011
rect 30607 14977 30616 15011
rect 30564 14968 30616 14977
rect 31024 14968 31076 15020
rect 33232 14968 33284 15020
rect 33876 14968 33928 15020
rect 46848 14968 46900 15020
rect 15752 14832 15804 14884
rect 18236 14832 18288 14884
rect 24768 14832 24820 14884
rect 23388 14764 23440 14816
rect 23480 14807 23532 14816
rect 23480 14773 23489 14807
rect 23489 14773 23523 14807
rect 23523 14773 23532 14807
rect 23480 14764 23532 14773
rect 23664 14764 23716 14816
rect 23848 14764 23900 14816
rect 26884 14832 26936 14884
rect 25044 14764 25096 14816
rect 29368 14764 29420 14816
rect 29460 14764 29512 14816
rect 30288 14832 30340 14884
rect 32404 14900 32456 14952
rect 32496 14832 32548 14884
rect 47768 14807 47820 14816
rect 47768 14773 47777 14807
rect 47777 14773 47811 14807
rect 47811 14773 47820 14807
rect 47768 14764 47820 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 19340 14560 19392 14612
rect 20260 14560 20312 14612
rect 21456 14492 21508 14544
rect 21732 14492 21784 14544
rect 1768 14356 1820 14408
rect 18696 14356 18748 14408
rect 20812 14356 20864 14408
rect 22836 14399 22888 14408
rect 22836 14365 22845 14399
rect 22845 14365 22879 14399
rect 22879 14365 22888 14399
rect 22836 14356 22888 14365
rect 23480 14560 23532 14612
rect 24492 14560 24544 14612
rect 26424 14560 26476 14612
rect 29552 14560 29604 14612
rect 30840 14560 30892 14612
rect 31944 14560 31996 14612
rect 32496 14560 32548 14612
rect 48044 14560 48096 14612
rect 24768 14492 24820 14544
rect 29368 14492 29420 14544
rect 31024 14492 31076 14544
rect 25044 14424 25096 14476
rect 27988 14356 28040 14408
rect 29276 14356 29328 14408
rect 32128 14424 32180 14476
rect 33324 14467 33376 14476
rect 33324 14433 33333 14467
rect 33333 14433 33367 14467
rect 33367 14433 33376 14467
rect 33324 14424 33376 14433
rect 24676 14288 24728 14340
rect 24860 14288 24912 14340
rect 27804 14331 27856 14340
rect 27804 14297 27813 14331
rect 27813 14297 27847 14331
rect 27847 14297 27856 14331
rect 27804 14288 27856 14297
rect 21180 14220 21232 14272
rect 24492 14220 24544 14272
rect 26148 14220 26200 14272
rect 27436 14220 27488 14272
rect 30564 14356 30616 14408
rect 30840 14399 30892 14408
rect 30840 14365 30849 14399
rect 30849 14365 30883 14399
rect 30883 14365 30892 14399
rect 30840 14356 30892 14365
rect 31392 14356 31444 14408
rect 31852 14399 31904 14408
rect 31852 14365 31861 14399
rect 31861 14365 31895 14399
rect 31895 14365 31904 14399
rect 31852 14356 31904 14365
rect 32036 14399 32088 14408
rect 32036 14365 32045 14399
rect 32045 14365 32079 14399
rect 32079 14365 32088 14399
rect 32036 14356 32088 14365
rect 32220 14399 32272 14408
rect 32220 14365 32229 14399
rect 32229 14365 32263 14399
rect 32263 14365 32272 14399
rect 32220 14356 32272 14365
rect 32312 14356 32364 14408
rect 47768 14424 47820 14476
rect 30656 14288 30708 14340
rect 30104 14220 30156 14272
rect 33232 14331 33284 14340
rect 33232 14297 33241 14331
rect 33241 14297 33275 14331
rect 33275 14297 33284 14331
rect 33232 14288 33284 14297
rect 46848 14288 46900 14340
rect 48136 14331 48188 14340
rect 48136 14297 48145 14331
rect 48145 14297 48179 14331
rect 48179 14297 48188 14331
rect 48136 14288 48188 14297
rect 32680 14220 32732 14272
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 17040 13880 17092 13932
rect 20168 14016 20220 14068
rect 27436 14016 27488 14068
rect 1952 13855 2004 13864
rect 1952 13821 1961 13855
rect 1961 13821 1995 13855
rect 1995 13821 2004 13855
rect 1952 13812 2004 13821
rect 2780 13855 2832 13864
rect 2780 13821 2789 13855
rect 2789 13821 2823 13855
rect 2823 13821 2832 13855
rect 17316 13855 17368 13864
rect 2780 13812 2832 13821
rect 17316 13821 17325 13855
rect 17325 13821 17359 13855
rect 17359 13821 17368 13855
rect 17316 13812 17368 13821
rect 18052 13855 18104 13864
rect 18052 13821 18061 13855
rect 18061 13821 18095 13855
rect 18095 13821 18104 13855
rect 18052 13812 18104 13821
rect 19432 13812 19484 13864
rect 20260 13812 20312 13864
rect 20720 13880 20772 13932
rect 23848 13948 23900 14000
rect 24492 13948 24544 14000
rect 26148 13948 26200 14000
rect 26884 13948 26936 14000
rect 29184 14016 29236 14068
rect 30932 14016 30984 14068
rect 31392 14059 31444 14068
rect 31392 14025 31401 14059
rect 31401 14025 31435 14059
rect 31435 14025 31444 14059
rect 31392 14016 31444 14025
rect 32128 14016 32180 14068
rect 46848 14059 46900 14068
rect 46848 14025 46857 14059
rect 46857 14025 46891 14059
rect 46891 14025 46900 14059
rect 46848 14016 46900 14025
rect 48044 14059 48096 14068
rect 48044 14025 48053 14059
rect 48053 14025 48087 14059
rect 48087 14025 48096 14059
rect 48044 14016 48096 14025
rect 32312 13948 32364 14000
rect 32680 13991 32732 14000
rect 32680 13957 32714 13991
rect 32714 13957 32732 13991
rect 32680 13948 32732 13957
rect 20996 13812 21048 13864
rect 23664 13812 23716 13864
rect 19524 13676 19576 13728
rect 23296 13719 23348 13728
rect 23296 13685 23305 13719
rect 23305 13685 23339 13719
rect 23339 13685 23348 13719
rect 23296 13676 23348 13685
rect 24124 13812 24176 13864
rect 27252 13880 27304 13932
rect 27896 13880 27948 13932
rect 29460 13923 29512 13932
rect 29460 13889 29469 13923
rect 29469 13889 29503 13923
rect 29503 13889 29512 13923
rect 29460 13880 29512 13889
rect 29644 13923 29696 13932
rect 29644 13889 29653 13923
rect 29653 13889 29687 13923
rect 29687 13889 29696 13923
rect 29644 13880 29696 13889
rect 31024 13923 31076 13932
rect 31024 13889 31033 13923
rect 31033 13889 31067 13923
rect 31067 13889 31076 13923
rect 31024 13880 31076 13889
rect 32404 13923 32456 13932
rect 24032 13744 24084 13796
rect 26424 13812 26476 13864
rect 26332 13744 26384 13796
rect 30656 13812 30708 13864
rect 30932 13812 30984 13864
rect 30012 13744 30064 13796
rect 30748 13744 30800 13796
rect 32404 13889 32413 13923
rect 32413 13889 32447 13923
rect 32447 13889 32456 13923
rect 32404 13880 32456 13889
rect 33784 13880 33836 13932
rect 47860 13923 47912 13932
rect 47860 13889 47869 13923
rect 47869 13889 47903 13923
rect 47903 13889 47912 13923
rect 47860 13880 47912 13889
rect 24584 13719 24636 13728
rect 24584 13685 24593 13719
rect 24593 13685 24627 13719
rect 24627 13685 24636 13719
rect 24584 13676 24636 13685
rect 24676 13676 24728 13728
rect 30840 13676 30892 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 1952 13472 2004 13524
rect 17316 13515 17368 13524
rect 17316 13481 17325 13515
rect 17325 13481 17359 13515
rect 17359 13481 17368 13515
rect 17316 13472 17368 13481
rect 1952 13268 2004 13320
rect 2320 13268 2372 13320
rect 7104 13268 7156 13320
rect 16856 13268 16908 13320
rect 21824 13472 21876 13524
rect 23848 13472 23900 13524
rect 24308 13472 24360 13524
rect 27252 13472 27304 13524
rect 29368 13472 29420 13524
rect 31024 13472 31076 13524
rect 19248 13379 19300 13388
rect 19248 13345 19257 13379
rect 19257 13345 19291 13379
rect 19291 13345 19300 13379
rect 19248 13336 19300 13345
rect 19524 13311 19576 13320
rect 19524 13277 19558 13311
rect 19558 13277 19576 13311
rect 19524 13268 19576 13277
rect 21364 13268 21416 13320
rect 23296 13268 23348 13320
rect 20168 13200 20220 13252
rect 25964 13404 26016 13456
rect 26240 13447 26292 13456
rect 26240 13413 26249 13447
rect 26249 13413 26283 13447
rect 26283 13413 26292 13447
rect 26240 13404 26292 13413
rect 29460 13404 29512 13456
rect 23480 13336 23532 13388
rect 24492 13336 24544 13388
rect 24768 13379 24820 13388
rect 24768 13345 24777 13379
rect 24777 13345 24811 13379
rect 24811 13345 24820 13379
rect 25504 13379 25556 13388
rect 24768 13336 24820 13345
rect 24676 13268 24728 13320
rect 25504 13345 25513 13379
rect 25513 13345 25547 13379
rect 25547 13345 25556 13379
rect 25504 13336 25556 13345
rect 27160 13336 27212 13388
rect 28172 13336 28224 13388
rect 32128 13379 32180 13388
rect 32128 13345 32137 13379
rect 32137 13345 32171 13379
rect 32171 13345 32180 13379
rect 32128 13336 32180 13345
rect 32312 13379 32364 13388
rect 32312 13345 32321 13379
rect 32321 13345 32355 13379
rect 32355 13345 32364 13379
rect 32312 13336 32364 13345
rect 25320 13311 25372 13320
rect 25320 13277 25329 13311
rect 25329 13277 25363 13311
rect 25363 13277 25372 13311
rect 25320 13268 25372 13277
rect 27804 13268 27856 13320
rect 27896 13311 27948 13320
rect 27896 13277 27905 13311
rect 27905 13277 27939 13311
rect 27939 13277 27948 13311
rect 27896 13268 27948 13277
rect 29276 13268 29328 13320
rect 30656 13311 30708 13320
rect 19156 13132 19208 13184
rect 20260 13132 20312 13184
rect 23388 13132 23440 13184
rect 24124 13132 24176 13184
rect 24952 13132 25004 13184
rect 27252 13132 27304 13184
rect 27896 13132 27948 13184
rect 29644 13132 29696 13184
rect 30656 13277 30665 13311
rect 30665 13277 30699 13311
rect 30699 13277 30708 13311
rect 30656 13268 30708 13277
rect 32220 13268 32272 13320
rect 30564 13132 30616 13184
rect 31116 13132 31168 13184
rect 32312 13132 32364 13184
rect 32772 13132 32824 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 3516 12792 3568 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 18236 12835 18288 12844
rect 18236 12801 18245 12835
rect 18245 12801 18279 12835
rect 18279 12801 18288 12835
rect 18236 12792 18288 12801
rect 19248 12792 19300 12844
rect 21272 12792 21324 12844
rect 23480 12928 23532 12980
rect 24768 12928 24820 12980
rect 27160 12971 27212 12980
rect 27160 12937 27169 12971
rect 27169 12937 27203 12971
rect 27203 12937 27212 12971
rect 27160 12928 27212 12937
rect 25596 12860 25648 12912
rect 27620 12860 27672 12912
rect 27804 12860 27856 12912
rect 30656 12860 30708 12912
rect 23204 12835 23256 12844
rect 1400 12767 1452 12776
rect 1400 12733 1409 12767
rect 1409 12733 1443 12767
rect 1443 12733 1452 12767
rect 1400 12724 1452 12733
rect 15844 12724 15896 12776
rect 20260 12724 20312 12776
rect 20168 12656 20220 12708
rect 23204 12801 23213 12835
rect 23213 12801 23247 12835
rect 23247 12801 23256 12835
rect 23204 12792 23256 12801
rect 23296 12792 23348 12844
rect 24032 12835 24084 12844
rect 24032 12801 24041 12835
rect 24041 12801 24075 12835
rect 24075 12801 24084 12835
rect 24032 12792 24084 12801
rect 24400 12792 24452 12844
rect 25320 12835 25372 12844
rect 25320 12801 25329 12835
rect 25329 12801 25363 12835
rect 25363 12801 25372 12835
rect 25320 12792 25372 12801
rect 23848 12724 23900 12776
rect 24124 12767 24176 12776
rect 24124 12733 24133 12767
rect 24133 12733 24167 12767
rect 24167 12733 24176 12767
rect 24124 12724 24176 12733
rect 24492 12724 24544 12776
rect 23480 12656 23532 12708
rect 16948 12631 17000 12640
rect 16948 12597 16957 12631
rect 16957 12597 16991 12631
rect 16991 12597 17000 12631
rect 16948 12588 17000 12597
rect 20720 12588 20772 12640
rect 22652 12631 22704 12640
rect 22652 12597 22661 12631
rect 22661 12597 22695 12631
rect 22695 12597 22704 12631
rect 22652 12588 22704 12597
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 24676 12588 24728 12640
rect 26240 12835 26292 12844
rect 26240 12801 26254 12835
rect 26254 12801 26288 12835
rect 26288 12801 26292 12835
rect 26240 12792 26292 12801
rect 27252 12835 27304 12844
rect 27252 12801 27261 12835
rect 27261 12801 27295 12835
rect 27295 12801 27304 12835
rect 29644 12835 29696 12844
rect 27252 12792 27304 12801
rect 29644 12801 29653 12835
rect 29653 12801 29687 12835
rect 29687 12801 29696 12835
rect 29644 12792 29696 12801
rect 29828 12835 29880 12844
rect 29828 12801 29837 12835
rect 29837 12801 29871 12835
rect 29871 12801 29880 12835
rect 29828 12792 29880 12801
rect 26332 12724 26384 12776
rect 26148 12656 26200 12708
rect 29736 12724 29788 12776
rect 30196 12792 30248 12844
rect 26424 12631 26476 12640
rect 26424 12597 26433 12631
rect 26433 12597 26467 12631
rect 26467 12597 26476 12631
rect 26424 12588 26476 12597
rect 26884 12588 26936 12640
rect 27160 12588 27212 12640
rect 30748 12656 30800 12708
rect 36636 12724 36688 12776
rect 46848 12724 46900 12776
rect 37832 12656 37884 12708
rect 30840 12588 30892 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 21272 12384 21324 12436
rect 24676 12427 24728 12436
rect 24676 12393 24685 12427
rect 24685 12393 24719 12427
rect 24719 12393 24728 12427
rect 24676 12384 24728 12393
rect 28080 12384 28132 12436
rect 29828 12384 29880 12436
rect 36452 12384 36504 12436
rect 45560 12384 45612 12436
rect 24584 12316 24636 12368
rect 22652 12248 22704 12300
rect 25044 12316 25096 12368
rect 27252 12316 27304 12368
rect 25320 12248 25372 12300
rect 19340 12180 19392 12232
rect 21364 12180 21416 12232
rect 23664 12223 23716 12232
rect 23664 12189 23673 12223
rect 23673 12189 23707 12223
rect 23707 12189 23716 12223
rect 23664 12180 23716 12189
rect 24032 12180 24084 12232
rect 24952 12223 25004 12232
rect 24952 12189 24961 12223
rect 24961 12189 24995 12223
rect 24995 12189 25004 12223
rect 24952 12180 25004 12189
rect 27528 12180 27580 12232
rect 28172 12180 28224 12232
rect 29644 12248 29696 12300
rect 20168 12112 20220 12164
rect 24860 12112 24912 12164
rect 26424 12155 26476 12164
rect 26424 12121 26458 12155
rect 26458 12121 26476 12155
rect 28080 12155 28132 12164
rect 26424 12112 26476 12121
rect 28080 12121 28089 12155
rect 28089 12121 28123 12155
rect 28123 12121 28132 12155
rect 28080 12112 28132 12121
rect 29552 12112 29604 12164
rect 29828 12223 29880 12232
rect 29828 12189 29837 12223
rect 29837 12189 29871 12223
rect 29871 12189 29880 12223
rect 30012 12223 30064 12232
rect 29828 12180 29880 12189
rect 30012 12189 30021 12223
rect 30021 12189 30055 12223
rect 30055 12189 30064 12223
rect 30012 12180 30064 12189
rect 30748 12112 30800 12164
rect 22100 12044 22152 12096
rect 22836 12087 22888 12096
rect 22836 12053 22845 12087
rect 22845 12053 22879 12087
rect 22879 12053 22888 12087
rect 22836 12044 22888 12053
rect 23388 12044 23440 12096
rect 25596 12044 25648 12096
rect 26056 12044 26108 12096
rect 26148 12044 26200 12096
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 20168 11883 20220 11892
rect 20168 11849 20177 11883
rect 20177 11849 20211 11883
rect 20211 11849 20220 11883
rect 20168 11840 20220 11849
rect 20444 11840 20496 11892
rect 20628 11840 20680 11892
rect 20812 11840 20864 11892
rect 21088 11840 21140 11892
rect 23480 11840 23532 11892
rect 25320 11840 25372 11892
rect 26056 11883 26108 11892
rect 26056 11849 26065 11883
rect 26065 11849 26099 11883
rect 26099 11849 26108 11883
rect 26056 11840 26108 11849
rect 26792 11840 26844 11892
rect 27344 11840 27396 11892
rect 27988 11840 28040 11892
rect 29460 11883 29512 11892
rect 29460 11849 29469 11883
rect 29469 11849 29503 11883
rect 29503 11849 29512 11883
rect 29460 11840 29512 11849
rect 16948 11815 17000 11824
rect 16948 11781 16957 11815
rect 16957 11781 16991 11815
rect 16991 11781 17000 11815
rect 16948 11772 17000 11781
rect 2228 11747 2280 11756
rect 2228 11713 2237 11747
rect 2237 11713 2271 11747
rect 2271 11713 2280 11747
rect 2228 11704 2280 11713
rect 11520 11704 11572 11756
rect 16764 11679 16816 11688
rect 16764 11645 16773 11679
rect 16773 11645 16807 11679
rect 16807 11645 16816 11679
rect 16764 11636 16816 11645
rect 18144 11679 18196 11688
rect 18144 11645 18153 11679
rect 18153 11645 18187 11679
rect 18187 11645 18196 11679
rect 18144 11636 18196 11645
rect 19616 11704 19668 11756
rect 20168 11704 20220 11756
rect 20260 11636 20312 11688
rect 20720 11704 20772 11756
rect 21272 11772 21324 11824
rect 22100 11747 22152 11756
rect 22100 11713 22109 11747
rect 22109 11713 22143 11747
rect 22143 11713 22152 11747
rect 22100 11704 22152 11713
rect 1584 11500 1636 11552
rect 2964 11543 3016 11552
rect 2964 11509 2973 11543
rect 2973 11509 3007 11543
rect 3007 11509 3016 11543
rect 2964 11500 3016 11509
rect 19064 11543 19116 11552
rect 19064 11509 19073 11543
rect 19073 11509 19107 11543
rect 19107 11509 19116 11543
rect 19064 11500 19116 11509
rect 20168 11568 20220 11620
rect 23204 11704 23256 11756
rect 25044 11704 25096 11756
rect 25780 11704 25832 11756
rect 27068 11704 27120 11756
rect 27620 11704 27672 11756
rect 22836 11636 22888 11688
rect 24492 11636 24544 11688
rect 24676 11636 24728 11688
rect 25596 11636 25648 11688
rect 26148 11679 26200 11688
rect 26148 11645 26157 11679
rect 26157 11645 26191 11679
rect 26191 11645 26200 11679
rect 26148 11636 26200 11645
rect 26332 11679 26384 11688
rect 26332 11645 26341 11679
rect 26341 11645 26375 11679
rect 26375 11645 26384 11679
rect 26332 11636 26384 11645
rect 29276 11747 29328 11756
rect 29276 11713 29285 11747
rect 29285 11713 29319 11747
rect 29319 11713 29328 11747
rect 29276 11704 29328 11713
rect 30472 11704 30524 11756
rect 36636 11704 36688 11756
rect 24860 11568 24912 11620
rect 25504 11568 25556 11620
rect 28632 11568 28684 11620
rect 29644 11636 29696 11688
rect 30656 11679 30708 11688
rect 21548 11500 21600 11552
rect 21916 11543 21968 11552
rect 21916 11509 21925 11543
rect 21925 11509 21959 11543
rect 21959 11509 21968 11543
rect 21916 11500 21968 11509
rect 28908 11500 28960 11552
rect 29552 11568 29604 11620
rect 30656 11645 30665 11679
rect 30665 11645 30699 11679
rect 30699 11645 30708 11679
rect 30656 11636 30708 11645
rect 30104 11568 30156 11620
rect 32496 11636 32548 11688
rect 46296 11500 46348 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 16764 11296 16816 11348
rect 19616 11339 19668 11348
rect 2964 11160 3016 11212
rect 3056 11203 3108 11212
rect 3056 11169 3065 11203
rect 3065 11169 3099 11203
rect 3099 11169 3108 11203
rect 19616 11305 19625 11339
rect 19625 11305 19659 11339
rect 19659 11305 19668 11339
rect 19616 11296 19668 11305
rect 22836 11296 22888 11348
rect 25596 11296 25648 11348
rect 25688 11296 25740 11348
rect 26240 11296 26292 11348
rect 27344 11296 27396 11348
rect 29276 11296 29328 11348
rect 30656 11296 30708 11348
rect 3056 11160 3108 11169
rect 17316 11135 17368 11144
rect 17316 11101 17325 11135
rect 17325 11101 17359 11135
rect 17359 11101 17368 11135
rect 17316 11092 17368 11101
rect 19064 11092 19116 11144
rect 19248 11135 19300 11144
rect 19248 11101 19257 11135
rect 19257 11101 19291 11135
rect 19291 11101 19300 11135
rect 19248 11092 19300 11101
rect 21088 11092 21140 11144
rect 21364 11135 21416 11144
rect 21364 11101 21373 11135
rect 21373 11101 21407 11135
rect 21407 11101 21416 11135
rect 21364 11092 21416 11101
rect 21916 11092 21968 11144
rect 24124 11092 24176 11144
rect 27160 11228 27212 11280
rect 27528 11228 27580 11280
rect 26332 11160 26384 11212
rect 27620 11135 27672 11144
rect 27620 11101 27629 11135
rect 27629 11101 27663 11135
rect 27663 11101 27672 11135
rect 27620 11092 27672 11101
rect 28080 11092 28132 11144
rect 28632 11135 28684 11144
rect 28632 11101 28641 11135
rect 28641 11101 28675 11135
rect 28675 11101 28684 11135
rect 28632 11092 28684 11101
rect 2872 11024 2924 11076
rect 19524 11024 19576 11076
rect 20444 11024 20496 11076
rect 24400 11067 24452 11076
rect 24400 11033 24409 11067
rect 24409 11033 24443 11067
rect 24443 11033 24452 11067
rect 24400 11024 24452 11033
rect 27528 11024 27580 11076
rect 30104 11203 30156 11212
rect 30104 11169 30113 11203
rect 30113 11169 30147 11203
rect 30147 11169 30156 11203
rect 30104 11160 30156 11169
rect 30748 11203 30800 11212
rect 30748 11169 30757 11203
rect 30757 11169 30791 11203
rect 30791 11169 30800 11203
rect 30748 11160 30800 11169
rect 46296 11203 46348 11212
rect 46296 11169 46305 11203
rect 46305 11169 46339 11203
rect 46339 11169 46348 11203
rect 46296 11160 46348 11169
rect 29920 11135 29972 11144
rect 29920 11101 29929 11135
rect 29929 11101 29963 11135
rect 29963 11101 29972 11135
rect 29920 11092 29972 11101
rect 30288 11092 30340 11144
rect 30840 11092 30892 11144
rect 46940 11024 46992 11076
rect 48136 11067 48188 11076
rect 48136 11033 48145 11067
rect 48145 11033 48179 11067
rect 48179 11033 48188 11067
rect 48136 11024 48188 11033
rect 19984 10956 20036 11008
rect 21272 10956 21324 11008
rect 27988 10999 28040 11008
rect 27988 10965 27997 10999
rect 27997 10965 28031 10999
rect 28031 10965 28040 10999
rect 27988 10956 28040 10965
rect 28448 10999 28500 11008
rect 28448 10965 28457 10999
rect 28457 10965 28491 10999
rect 28491 10965 28500 10999
rect 28448 10956 28500 10965
rect 29552 10999 29604 11008
rect 29552 10965 29561 10999
rect 29561 10965 29595 10999
rect 29595 10965 29604 10999
rect 29552 10956 29604 10965
rect 30012 10999 30064 11008
rect 30012 10965 30021 10999
rect 30021 10965 30055 10999
rect 30055 10965 30064 10999
rect 30012 10956 30064 10965
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 27528 10752 27580 10804
rect 29368 10752 29420 10804
rect 46940 10795 46992 10804
rect 46940 10761 46949 10795
rect 46949 10761 46983 10795
rect 46983 10761 46992 10795
rect 46940 10752 46992 10761
rect 20260 10684 20312 10736
rect 27160 10727 27212 10736
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 14556 10616 14608 10668
rect 19156 10616 19208 10668
rect 19616 10616 19668 10668
rect 20628 10616 20680 10668
rect 24032 10659 24084 10668
rect 24032 10625 24041 10659
rect 24041 10625 24075 10659
rect 24075 10625 24084 10659
rect 24032 10616 24084 10625
rect 27160 10693 27169 10727
rect 27169 10693 27203 10727
rect 27203 10693 27212 10727
rect 27160 10684 27212 10693
rect 26240 10659 26292 10668
rect 26240 10625 26249 10659
rect 26249 10625 26283 10659
rect 26283 10625 26292 10659
rect 26240 10616 26292 10625
rect 2872 10591 2924 10600
rect 2872 10557 2881 10591
rect 2881 10557 2915 10591
rect 2915 10557 2924 10591
rect 2872 10548 2924 10557
rect 23112 10548 23164 10600
rect 26332 10548 26384 10600
rect 27344 10616 27396 10668
rect 27712 10684 27764 10736
rect 28908 10684 28960 10736
rect 29276 10616 29328 10668
rect 29460 10684 29512 10736
rect 29736 10659 29788 10668
rect 29736 10625 29745 10659
rect 29745 10625 29779 10659
rect 29779 10625 29788 10659
rect 29736 10616 29788 10625
rect 30288 10659 30340 10668
rect 30288 10625 30297 10659
rect 30297 10625 30331 10659
rect 30331 10625 30340 10659
rect 30288 10616 30340 10625
rect 30564 10616 30616 10668
rect 30932 10616 30984 10668
rect 46848 10659 46900 10668
rect 46848 10625 46857 10659
rect 46857 10625 46891 10659
rect 46891 10625 46900 10659
rect 46848 10616 46900 10625
rect 47768 10659 47820 10668
rect 47768 10625 47777 10659
rect 47777 10625 47811 10659
rect 47811 10625 47820 10659
rect 47768 10616 47820 10625
rect 30012 10591 30064 10600
rect 23480 10480 23532 10532
rect 24584 10480 24636 10532
rect 3516 10455 3568 10464
rect 3516 10421 3525 10455
rect 3525 10421 3559 10455
rect 3559 10421 3568 10455
rect 3516 10412 3568 10421
rect 19064 10455 19116 10464
rect 19064 10421 19073 10455
rect 19073 10421 19107 10455
rect 19107 10421 19116 10455
rect 19064 10412 19116 10421
rect 27068 10480 27120 10532
rect 30012 10557 30021 10591
rect 30021 10557 30055 10591
rect 30055 10557 30064 10591
rect 30012 10548 30064 10557
rect 30104 10591 30156 10600
rect 30104 10557 30113 10591
rect 30113 10557 30147 10591
rect 30147 10557 30156 10591
rect 30104 10548 30156 10557
rect 26332 10455 26384 10464
rect 26332 10421 26341 10455
rect 26341 10421 26375 10455
rect 26375 10421 26384 10455
rect 26332 10412 26384 10421
rect 26516 10412 26568 10464
rect 27344 10412 27396 10464
rect 30656 10480 30708 10532
rect 30932 10480 30984 10532
rect 29368 10412 29420 10464
rect 30840 10412 30892 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 19616 10251 19668 10260
rect 19616 10217 19625 10251
rect 19625 10217 19659 10251
rect 19659 10217 19668 10251
rect 19616 10208 19668 10217
rect 21548 10208 21600 10260
rect 20628 10140 20680 10192
rect 3516 10072 3568 10124
rect 20260 10072 20312 10124
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 1584 9979 1636 9988
rect 1584 9945 1593 9979
rect 1593 9945 1627 9979
rect 1627 9945 1636 9979
rect 1584 9936 1636 9945
rect 3240 9979 3292 9988
rect 3240 9945 3249 9979
rect 3249 9945 3283 9979
rect 3283 9945 3292 9979
rect 3240 9936 3292 9945
rect 19340 9936 19392 9988
rect 20720 10047 20772 10056
rect 20720 10013 20729 10047
rect 20729 10013 20763 10047
rect 20763 10013 20772 10047
rect 20720 10004 20772 10013
rect 23112 10047 23164 10056
rect 23112 10013 23121 10047
rect 23121 10013 23155 10047
rect 23155 10013 23164 10047
rect 23480 10208 23532 10260
rect 24032 10208 24084 10260
rect 26240 10208 26292 10260
rect 26424 10208 26476 10260
rect 24676 10140 24728 10192
rect 24400 10072 24452 10124
rect 26516 10115 26568 10124
rect 26516 10081 26525 10115
rect 26525 10081 26559 10115
rect 26559 10081 26568 10115
rect 26516 10072 26568 10081
rect 27896 10140 27948 10192
rect 28540 10140 28592 10192
rect 29828 10208 29880 10260
rect 30012 10208 30064 10260
rect 30564 10140 30616 10192
rect 28448 10072 28500 10124
rect 23112 10004 23164 10013
rect 23480 10047 23532 10056
rect 23480 10013 23489 10047
rect 23489 10013 23523 10047
rect 23523 10013 23532 10047
rect 23480 10004 23532 10013
rect 27988 10004 28040 10056
rect 20904 9868 20956 9920
rect 22192 9868 22244 9920
rect 23296 9868 23348 9920
rect 23480 9868 23532 9920
rect 25136 9936 25188 9988
rect 26056 9936 26108 9988
rect 28908 10004 28960 10056
rect 29552 10047 29604 10056
rect 29552 10013 29561 10047
rect 29561 10013 29595 10047
rect 29595 10013 29604 10047
rect 29552 10004 29604 10013
rect 23848 9911 23900 9920
rect 23848 9877 23857 9911
rect 23857 9877 23891 9911
rect 23891 9877 23900 9911
rect 23848 9868 23900 9877
rect 24584 9868 24636 9920
rect 25780 9868 25832 9920
rect 26424 9911 26476 9920
rect 26424 9877 26433 9911
rect 26433 9877 26467 9911
rect 26467 9877 26476 9911
rect 26424 9868 26476 9877
rect 28172 9868 28224 9920
rect 30656 10004 30708 10056
rect 30840 10047 30892 10056
rect 30840 10013 30874 10047
rect 30874 10013 30892 10047
rect 30840 10004 30892 10013
rect 42432 9936 42484 9988
rect 46848 9936 46900 9988
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 2964 9596 3016 9648
rect 18052 9664 18104 9716
rect 20720 9664 20772 9716
rect 24400 9664 24452 9716
rect 28264 9664 28316 9716
rect 29460 9664 29512 9716
rect 29736 9664 29788 9716
rect 17316 9528 17368 9580
rect 21088 9596 21140 9648
rect 19064 9528 19116 9580
rect 19248 9528 19300 9580
rect 21916 9528 21968 9580
rect 25964 9596 26016 9648
rect 23848 9528 23900 9580
rect 25780 9528 25832 9580
rect 26516 9596 26568 9648
rect 26424 9528 26476 9580
rect 28632 9528 28684 9580
rect 29000 9528 29052 9580
rect 29828 9528 29880 9580
rect 26056 9503 26108 9512
rect 26056 9469 26065 9503
rect 26065 9469 26099 9503
rect 26099 9469 26108 9503
rect 28448 9503 28500 9512
rect 26056 9460 26108 9469
rect 28448 9469 28457 9503
rect 28457 9469 28491 9503
rect 28491 9469 28500 9503
rect 28448 9460 28500 9469
rect 28540 9503 28592 9512
rect 28540 9469 28549 9503
rect 28549 9469 28583 9503
rect 28583 9469 28592 9503
rect 28540 9460 28592 9469
rect 26332 9392 26384 9444
rect 27620 9392 27672 9444
rect 19340 9324 19392 9376
rect 26240 9324 26292 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 17316 9027 17368 9036
rect 17316 8993 17325 9027
rect 17325 8993 17359 9027
rect 17359 8993 17368 9027
rect 17316 8984 17368 8993
rect 20260 9120 20312 9172
rect 25780 9120 25832 9172
rect 27344 9163 27396 9172
rect 19984 9052 20036 9104
rect 25964 9027 26016 9036
rect 25964 8993 25973 9027
rect 25973 8993 26007 9027
rect 26007 8993 26016 9027
rect 25964 8984 26016 8993
rect 27344 9129 27353 9163
rect 27353 9129 27387 9163
rect 27387 9129 27396 9163
rect 27344 9120 27396 9129
rect 27436 9120 27488 9172
rect 32588 9120 32640 9172
rect 28540 9052 28592 9104
rect 30104 9052 30156 9104
rect 28264 8984 28316 9036
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 20168 8959 20220 8968
rect 20168 8925 20177 8959
rect 20177 8925 20211 8959
rect 20211 8925 20220 8959
rect 20168 8916 20220 8925
rect 20720 8916 20772 8968
rect 20904 8959 20956 8968
rect 20904 8925 20938 8959
rect 20938 8925 20956 8959
rect 20904 8916 20956 8925
rect 26240 8959 26292 8968
rect 26240 8925 26274 8959
rect 26274 8925 26292 8959
rect 26240 8916 26292 8925
rect 28172 8959 28224 8968
rect 28172 8925 28181 8959
rect 28181 8925 28215 8959
rect 28215 8925 28224 8959
rect 28172 8916 28224 8925
rect 28448 9027 28500 9036
rect 28448 8993 28457 9027
rect 28457 8993 28491 9027
rect 28491 8993 28500 9027
rect 28448 8984 28500 8993
rect 29276 8984 29328 9036
rect 29736 8984 29788 9036
rect 28540 8959 28592 8968
rect 28540 8925 28549 8959
rect 28549 8925 28583 8959
rect 28583 8925 28592 8959
rect 28540 8916 28592 8925
rect 28632 8916 28684 8968
rect 20812 8848 20864 8900
rect 26884 8848 26936 8900
rect 28816 8848 28868 8900
rect 30748 8848 30800 8900
rect 47952 8891 48004 8900
rect 47952 8857 47961 8891
rect 47961 8857 47995 8891
rect 47995 8857 48004 8891
rect 47952 8848 48004 8857
rect 18880 8780 18932 8832
rect 20720 8780 20772 8832
rect 21088 8780 21140 8832
rect 21916 8780 21968 8832
rect 28908 8823 28960 8832
rect 28908 8789 28917 8823
rect 28917 8789 28951 8823
rect 28951 8789 28960 8823
rect 28908 8780 28960 8789
rect 38292 8780 38344 8832
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 27528 8576 27580 8628
rect 29736 8619 29788 8628
rect 1860 8483 1912 8492
rect 1860 8449 1869 8483
rect 1869 8449 1903 8483
rect 1903 8449 1912 8483
rect 1860 8440 1912 8449
rect 19340 8508 19392 8560
rect 18696 8415 18748 8424
rect 18696 8381 18705 8415
rect 18705 8381 18739 8415
rect 18739 8381 18748 8415
rect 18696 8372 18748 8381
rect 19432 8415 19484 8424
rect 19432 8381 19441 8415
rect 19441 8381 19475 8415
rect 19475 8381 19484 8415
rect 19432 8372 19484 8381
rect 20812 8372 20864 8424
rect 21824 8372 21876 8424
rect 26424 8372 26476 8424
rect 16672 8304 16724 8356
rect 20168 8304 20220 8356
rect 27436 8304 27488 8356
rect 28908 8440 28960 8492
rect 29736 8585 29745 8619
rect 29745 8585 29779 8619
rect 29779 8585 29788 8619
rect 29736 8576 29788 8585
rect 30748 8576 30800 8628
rect 30472 8483 30524 8492
rect 30472 8449 30481 8483
rect 30481 8449 30515 8483
rect 30515 8449 30524 8483
rect 30472 8440 30524 8449
rect 32588 8440 32640 8492
rect 47768 8483 47820 8492
rect 47768 8449 47777 8483
rect 47777 8449 47811 8483
rect 47811 8449 47820 8483
rect 47768 8440 47820 8449
rect 31852 8372 31904 8424
rect 30656 8304 30708 8356
rect 30196 8279 30248 8288
rect 30196 8245 30205 8279
rect 30205 8245 30239 8279
rect 30239 8245 30248 8279
rect 30196 8236 30248 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 18696 8032 18748 8084
rect 19984 8032 20036 8084
rect 20720 8032 20772 8084
rect 21732 8032 21784 8084
rect 23848 8032 23900 8084
rect 31852 8075 31904 8084
rect 21364 7964 21416 8016
rect 16488 7896 16540 7948
rect 1860 7803 1912 7812
rect 1860 7769 1869 7803
rect 1869 7769 1903 7803
rect 1903 7769 1912 7803
rect 1860 7760 1912 7769
rect 18880 7828 18932 7880
rect 19248 7760 19300 7812
rect 19340 7760 19392 7812
rect 21732 7828 21784 7880
rect 22100 7964 22152 8016
rect 22284 7964 22336 8016
rect 22192 7871 22244 7880
rect 22192 7837 22201 7871
rect 22201 7837 22235 7871
rect 22235 7837 22244 7871
rect 22192 7828 22244 7837
rect 22652 7828 22704 7880
rect 23664 7964 23716 8016
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 26884 7871 26936 7880
rect 26884 7837 26893 7871
rect 26893 7837 26927 7871
rect 26927 7837 26936 7871
rect 26884 7828 26936 7837
rect 22100 7760 22152 7812
rect 22284 7760 22336 7812
rect 27436 7828 27488 7880
rect 27528 7760 27580 7812
rect 30656 7828 30708 7880
rect 31852 8041 31861 8075
rect 31861 8041 31895 8075
rect 31895 8041 31904 8075
rect 31852 8032 31904 8041
rect 18972 7692 19024 7744
rect 20904 7735 20956 7744
rect 20904 7701 20913 7735
rect 20913 7701 20947 7735
rect 20947 7701 20956 7735
rect 20904 7692 20956 7701
rect 21456 7692 21508 7744
rect 24492 7692 24544 7744
rect 26608 7735 26660 7744
rect 26608 7701 26617 7735
rect 26617 7701 26651 7735
rect 26651 7701 26660 7735
rect 26608 7692 26660 7701
rect 26976 7692 27028 7744
rect 28264 7760 28316 7812
rect 30196 7760 30248 7812
rect 29644 7692 29696 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 22192 7488 22244 7540
rect 25228 7488 25280 7540
rect 19248 7420 19300 7472
rect 18880 7395 18932 7404
rect 18880 7361 18889 7395
rect 18889 7361 18923 7395
rect 18923 7361 18932 7395
rect 18880 7352 18932 7361
rect 20812 7352 20864 7404
rect 23756 7352 23808 7404
rect 26608 7420 26660 7472
rect 27804 7352 27856 7404
rect 29644 7395 29696 7404
rect 29644 7361 29653 7395
rect 29653 7361 29687 7395
rect 29687 7361 29696 7395
rect 29644 7352 29696 7361
rect 45744 7352 45796 7404
rect 19340 7284 19392 7336
rect 18696 7216 18748 7268
rect 21088 7284 21140 7336
rect 2044 7191 2096 7200
rect 2044 7157 2053 7191
rect 2053 7157 2087 7191
rect 2087 7157 2096 7191
rect 2044 7148 2096 7157
rect 25964 7284 26016 7336
rect 29828 7327 29880 7336
rect 29828 7293 29837 7327
rect 29837 7293 29871 7327
rect 29871 7293 29880 7327
rect 29828 7284 29880 7293
rect 29644 7216 29696 7268
rect 24952 7148 25004 7200
rect 25044 7191 25096 7200
rect 25044 7157 25053 7191
rect 25053 7157 25087 7191
rect 25087 7157 25096 7191
rect 25044 7148 25096 7157
rect 26700 7148 26752 7200
rect 28264 7148 28316 7200
rect 46480 7148 46532 7200
rect 47768 7191 47820 7200
rect 47768 7157 47777 7191
rect 47777 7157 47811 7191
rect 47811 7157 47820 7191
rect 47768 7148 47820 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 21824 6944 21876 6996
rect 22100 6944 22152 6996
rect 26884 6944 26936 6996
rect 29828 6987 29880 6996
rect 29828 6953 29837 6987
rect 29837 6953 29871 6987
rect 29871 6953 29880 6987
rect 29828 6944 29880 6953
rect 2044 6808 2096 6860
rect 2780 6851 2832 6860
rect 2780 6817 2789 6851
rect 2789 6817 2823 6851
rect 2823 6817 2832 6851
rect 2780 6808 2832 6817
rect 19340 6851 19392 6860
rect 19340 6817 19349 6851
rect 19349 6817 19383 6851
rect 19383 6817 19392 6851
rect 19340 6808 19392 6817
rect 20812 6808 20864 6860
rect 21088 6851 21140 6860
rect 21088 6817 21097 6851
rect 21097 6817 21131 6851
rect 21131 6817 21140 6851
rect 21088 6808 21140 6817
rect 23756 6808 23808 6860
rect 26700 6851 26752 6860
rect 26700 6817 26709 6851
rect 26709 6817 26743 6851
rect 26743 6817 26752 6851
rect 26700 6808 26752 6817
rect 26976 6851 27028 6860
rect 26976 6817 26985 6851
rect 26985 6817 27019 6851
rect 27019 6817 27028 6851
rect 26976 6808 27028 6817
rect 37096 6808 37148 6860
rect 45652 6808 45704 6860
rect 46480 6851 46532 6860
rect 46480 6817 46489 6851
rect 46489 6817 46523 6851
rect 46523 6817 46532 6851
rect 46480 6808 46532 6817
rect 48136 6851 48188 6860
rect 48136 6817 48145 6851
rect 48145 6817 48179 6851
rect 48179 6817 48188 6851
rect 48136 6808 48188 6817
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 2228 6672 2280 6724
rect 15200 6672 15252 6724
rect 20720 6740 20772 6792
rect 20904 6740 20956 6792
rect 23388 6740 23440 6792
rect 23572 6783 23624 6792
rect 23572 6749 23581 6783
rect 23581 6749 23615 6783
rect 23615 6749 23624 6783
rect 23572 6740 23624 6749
rect 23664 6783 23716 6792
rect 23664 6749 23673 6783
rect 23673 6749 23707 6783
rect 23707 6749 23716 6783
rect 23664 6740 23716 6749
rect 24032 6740 24084 6792
rect 24952 6740 25004 6792
rect 25964 6740 26016 6792
rect 21456 6672 21508 6724
rect 24492 6672 24544 6724
rect 27896 6740 27948 6792
rect 28264 6672 28316 6724
rect 37188 6672 37240 6724
rect 45560 6672 45612 6724
rect 47768 6672 47820 6724
rect 21548 6604 21600 6656
rect 23572 6604 23624 6656
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 2228 6443 2280 6452
rect 2228 6409 2237 6443
rect 2237 6409 2271 6443
rect 2271 6409 2280 6443
rect 2228 6400 2280 6409
rect 22192 6443 22244 6452
rect 22192 6409 22201 6443
rect 22201 6409 22235 6443
rect 22235 6409 22244 6443
rect 22192 6400 22244 6409
rect 23664 6400 23716 6452
rect 22100 6332 22152 6384
rect 25044 6332 25096 6384
rect 2136 6307 2188 6316
rect 2136 6273 2145 6307
rect 2145 6273 2179 6307
rect 2179 6273 2188 6307
rect 2136 6264 2188 6273
rect 22284 6196 22336 6248
rect 23388 6264 23440 6316
rect 38660 6400 38712 6452
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 3424 5856 3476 5908
rect 23480 5856 23532 5908
rect 25412 5856 25464 5908
rect 26976 5788 27028 5840
rect 2136 5652 2188 5704
rect 3056 5559 3108 5568
rect 3056 5525 3065 5559
rect 3065 5525 3099 5559
rect 3099 5525 3108 5559
rect 3056 5516 3108 5525
rect 25872 5652 25924 5704
rect 47400 5695 47452 5704
rect 47400 5661 47409 5695
rect 47409 5661 47443 5695
rect 47443 5661 47452 5695
rect 47400 5652 47452 5661
rect 35348 5584 35400 5636
rect 47952 5627 48004 5636
rect 47952 5593 47961 5627
rect 47961 5593 47995 5627
rect 47995 5593 48004 5627
rect 47952 5584 48004 5593
rect 26792 5516 26844 5568
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 3056 5244 3108 5296
rect 2136 5219 2188 5228
rect 2136 5185 2145 5219
rect 2145 5185 2179 5219
rect 2179 5185 2188 5219
rect 2136 5176 2188 5185
rect 46848 5219 46900 5228
rect 46848 5185 46857 5219
rect 46857 5185 46891 5219
rect 46891 5185 46900 5219
rect 46848 5176 46900 5185
rect 47492 5176 47544 5228
rect 47584 5219 47636 5228
rect 47584 5185 47593 5219
rect 47593 5185 47627 5219
rect 47627 5185 47636 5219
rect 47584 5176 47636 5185
rect 48228 5176 48280 5228
rect 2780 5151 2832 5160
rect 2780 5117 2789 5151
rect 2789 5117 2823 5151
rect 2823 5117 2832 5151
rect 2780 5108 2832 5117
rect 36360 5108 36412 5160
rect 47032 5108 47084 5160
rect 1400 4972 1452 5024
rect 46940 5015 46992 5024
rect 46940 4981 46949 5015
rect 46949 4981 46983 5015
rect 46983 4981 46992 5015
rect 46940 4972 46992 4981
rect 47676 5015 47728 5024
rect 47676 4981 47685 5015
rect 47685 4981 47719 5015
rect 47719 4981 47728 5015
rect 47676 4972 47728 4981
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 35440 4768 35492 4820
rect 45560 4768 45612 4820
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 21916 4632 21968 4684
rect 34796 4632 34848 4684
rect 37372 4632 37424 4684
rect 43076 4632 43128 4684
rect 43260 4675 43312 4684
rect 43260 4641 43269 4675
rect 43269 4641 43303 4675
rect 43303 4641 43312 4675
rect 43260 4632 43312 4641
rect 47400 4700 47452 4752
rect 47676 4632 47728 4684
rect 48136 4675 48188 4684
rect 48136 4641 48145 4675
rect 48145 4641 48179 4675
rect 48179 4641 48188 4675
rect 48136 4632 48188 4641
rect 3240 4607 3292 4616
rect 3240 4573 3249 4607
rect 3249 4573 3283 4607
rect 3283 4573 3292 4607
rect 3240 4564 3292 4573
rect 3792 4607 3844 4616
rect 3792 4573 3801 4607
rect 3801 4573 3835 4607
rect 3835 4573 3844 4607
rect 3792 4564 3844 4573
rect 6276 4607 6328 4616
rect 6276 4573 6285 4607
rect 6285 4573 6319 4607
rect 6319 4573 6328 4607
rect 6276 4564 6328 4573
rect 7196 4564 7248 4616
rect 8024 4607 8076 4616
rect 8024 4573 8033 4607
rect 8033 4573 8067 4607
rect 8067 4573 8076 4607
rect 8024 4564 8076 4573
rect 30472 4607 30524 4616
rect 30472 4573 30481 4607
rect 30481 4573 30515 4607
rect 30515 4573 30524 4607
rect 30472 4564 30524 4573
rect 30840 4564 30892 4616
rect 44732 4564 44784 4616
rect 45836 4607 45888 4616
rect 45836 4573 45845 4607
rect 45845 4573 45879 4607
rect 45879 4573 45888 4607
rect 45836 4564 45888 4573
rect 22192 4539 22244 4548
rect 22192 4505 22201 4539
rect 22201 4505 22235 4539
rect 22235 4505 22244 4539
rect 22192 4496 22244 4505
rect 34520 4496 34572 4548
rect 42064 4539 42116 4548
rect 42064 4505 42073 4539
rect 42073 4505 42107 4539
rect 42107 4505 42116 4539
rect 42064 4496 42116 4505
rect 8116 4471 8168 4480
rect 8116 4437 8125 4471
rect 8125 4437 8159 4471
rect 8159 4437 8168 4471
rect 8116 4428 8168 4437
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 22192 4224 22244 4276
rect 42064 4224 42116 4276
rect 3424 4156 3476 4208
rect 8116 4199 8168 4208
rect 1952 4088 2004 4140
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 6368 4131 6420 4140
rect 6368 4097 6377 4131
rect 6377 4097 6411 4131
rect 6411 4097 6420 4131
rect 6368 4088 6420 4097
rect 2136 4020 2188 4072
rect 6184 4020 6236 4072
rect 8116 4165 8125 4199
rect 8125 4165 8159 4199
rect 8159 4165 8168 4199
rect 8116 4156 8168 4165
rect 10232 4156 10284 4208
rect 17960 4156 18012 4208
rect 7012 4131 7064 4140
rect 7012 4097 7021 4131
rect 7021 4097 7055 4131
rect 7055 4097 7064 4131
rect 7932 4131 7984 4140
rect 7012 4088 7064 4097
rect 7932 4097 7941 4131
rect 7941 4097 7975 4131
rect 7975 4097 7984 4131
rect 7932 4088 7984 4097
rect 2504 3952 2556 4004
rect 12532 4131 12584 4140
rect 12532 4097 12541 4131
rect 12541 4097 12575 4131
rect 12575 4097 12584 4131
rect 12532 4088 12584 4097
rect 14924 4088 14976 4140
rect 22560 4131 22612 4140
rect 22560 4097 22569 4131
rect 22569 4097 22603 4131
rect 22603 4097 22612 4131
rect 29460 4156 29512 4208
rect 22560 4088 22612 4097
rect 30196 4088 30248 4140
rect 31300 4088 31352 4140
rect 1584 3927 1636 3936
rect 1584 3893 1593 3927
rect 1593 3893 1627 3927
rect 1627 3893 1636 3927
rect 1584 3884 1636 3893
rect 1676 3884 1728 3936
rect 2872 3884 2924 3936
rect 3516 3884 3568 3936
rect 5172 3884 5224 3936
rect 5540 3884 5592 3936
rect 7104 3927 7156 3936
rect 7104 3893 7113 3927
rect 7113 3893 7147 3927
rect 7147 3893 7156 3927
rect 7104 3884 7156 3893
rect 7932 3884 7984 3936
rect 10692 4020 10744 4072
rect 12440 4020 12492 4072
rect 13176 4063 13228 4072
rect 13176 4029 13185 4063
rect 13185 4029 13219 4063
rect 13219 4029 13228 4063
rect 13176 4020 13228 4029
rect 10324 3952 10376 4004
rect 12348 3952 12400 4004
rect 13544 4020 13596 4072
rect 17224 4020 17276 4072
rect 22468 4020 22520 4072
rect 26424 4020 26476 4072
rect 28356 4020 28408 4072
rect 11888 3884 11940 3936
rect 12532 3884 12584 3936
rect 24400 3952 24452 4004
rect 37832 4131 37884 4140
rect 37832 4097 37841 4131
rect 37841 4097 37875 4131
rect 37875 4097 37884 4131
rect 37832 4088 37884 4097
rect 42340 4088 42392 4140
rect 42432 4131 42484 4140
rect 42432 4097 42441 4131
rect 42441 4097 42475 4131
rect 42475 4097 42484 4131
rect 42432 4088 42484 4097
rect 46756 4156 46808 4208
rect 17316 3884 17368 3936
rect 20996 3927 21048 3936
rect 20996 3893 21005 3927
rect 21005 3893 21039 3927
rect 21039 3893 21048 3927
rect 20996 3884 21048 3893
rect 23388 3884 23440 3936
rect 25688 3884 25740 3936
rect 29736 3884 29788 3936
rect 31024 3884 31076 3936
rect 31484 3927 31536 3936
rect 31484 3893 31493 3927
rect 31493 3893 31527 3927
rect 31527 3893 31536 3927
rect 31484 3884 31536 3893
rect 32128 3884 32180 3936
rect 36268 3884 36320 3936
rect 38752 3884 38804 3936
rect 40776 3884 40828 3936
rect 42432 3884 42484 3936
rect 43996 4088 44048 4140
rect 45468 4088 45520 4140
rect 43812 4020 43864 4072
rect 44456 4020 44508 4072
rect 44824 3952 44876 4004
rect 46848 3952 46900 4004
rect 45744 3884 45796 3936
rect 46204 3884 46256 3936
rect 48044 3927 48096 3936
rect 48044 3893 48053 3927
rect 48053 3893 48087 3927
rect 48087 3893 48096 3927
rect 48044 3884 48096 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 2964 3680 3016 3732
rect 12440 3680 12492 3732
rect 1676 3544 1728 3596
rect 1860 3587 1912 3596
rect 1860 3553 1869 3587
rect 1869 3553 1903 3587
rect 1903 3553 1912 3587
rect 1860 3544 1912 3553
rect 3884 3476 3936 3528
rect 7932 3612 7984 3664
rect 8024 3612 8076 3664
rect 17224 3680 17276 3732
rect 17592 3680 17644 3732
rect 19432 3680 19484 3732
rect 22652 3723 22704 3732
rect 22652 3689 22661 3723
rect 22661 3689 22695 3723
rect 22695 3689 22704 3723
rect 22652 3680 22704 3689
rect 23296 3680 23348 3732
rect 33784 3680 33836 3732
rect 43076 3723 43128 3732
rect 43076 3689 43085 3723
rect 43085 3689 43119 3723
rect 43119 3689 43128 3723
rect 43076 3680 43128 3689
rect 43812 3723 43864 3732
rect 43812 3689 43821 3723
rect 43821 3689 43855 3723
rect 43855 3689 43864 3723
rect 43812 3680 43864 3689
rect 43996 3680 44048 3732
rect 47584 3680 47636 3732
rect 5172 3587 5224 3596
rect 5172 3553 5181 3587
rect 5181 3553 5215 3587
rect 5215 3553 5224 3587
rect 5172 3544 5224 3553
rect 5540 3544 5592 3596
rect 3976 3408 4028 3460
rect 3700 3340 3752 3392
rect 5172 3408 5224 3460
rect 7012 3544 7064 3596
rect 12808 3587 12860 3596
rect 12808 3553 12817 3587
rect 12817 3553 12851 3587
rect 12851 3553 12860 3587
rect 12808 3544 12860 3553
rect 9036 3476 9088 3528
rect 10508 3476 10560 3528
rect 11704 3519 11756 3528
rect 11704 3485 11713 3519
rect 11713 3485 11747 3519
rect 11747 3485 11756 3519
rect 11704 3476 11756 3485
rect 6920 3408 6972 3460
rect 11888 3451 11940 3460
rect 11888 3417 11897 3451
rect 11897 3417 11931 3451
rect 11931 3417 11940 3451
rect 11888 3408 11940 3417
rect 12440 3408 12492 3460
rect 18328 3544 18380 3596
rect 14924 3476 14976 3528
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 11520 3340 11572 3392
rect 11612 3340 11664 3392
rect 15476 3340 15528 3392
rect 17500 3340 17552 3392
rect 30012 3612 30064 3664
rect 30196 3612 30248 3664
rect 32404 3612 32456 3664
rect 35808 3612 35860 3664
rect 45468 3612 45520 3664
rect 20628 3544 20680 3596
rect 22468 3544 22520 3596
rect 25504 3544 25556 3596
rect 25688 3587 25740 3596
rect 25688 3553 25697 3587
rect 25697 3553 25731 3587
rect 25731 3553 25740 3587
rect 25688 3544 25740 3553
rect 26424 3587 26476 3596
rect 26424 3553 26433 3587
rect 26433 3553 26467 3587
rect 26467 3553 26476 3587
rect 26424 3544 26476 3553
rect 30840 3587 30892 3596
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 23204 3476 23256 3528
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 29552 3519 29604 3528
rect 23296 3476 23348 3485
rect 29552 3485 29561 3519
rect 29561 3485 29595 3519
rect 29595 3485 29604 3519
rect 29552 3476 29604 3485
rect 30196 3519 30248 3528
rect 30196 3485 30205 3519
rect 30205 3485 30239 3519
rect 30239 3485 30248 3519
rect 30196 3476 30248 3485
rect 23572 3340 23624 3392
rect 26148 3408 26200 3460
rect 30840 3553 30849 3587
rect 30849 3553 30883 3587
rect 30883 3553 30892 3587
rect 30840 3544 30892 3553
rect 31024 3587 31076 3596
rect 31024 3553 31033 3587
rect 31033 3553 31067 3587
rect 31067 3553 31076 3587
rect 31024 3544 31076 3553
rect 31576 3587 31628 3596
rect 31576 3553 31585 3587
rect 31585 3553 31619 3587
rect 31619 3553 31628 3587
rect 31576 3544 31628 3553
rect 36268 3587 36320 3596
rect 36268 3553 36277 3587
rect 36277 3553 36311 3587
rect 36311 3553 36320 3587
rect 36268 3544 36320 3553
rect 36728 3587 36780 3596
rect 36728 3553 36737 3587
rect 36737 3553 36771 3587
rect 36771 3553 36780 3587
rect 36728 3544 36780 3553
rect 40776 3587 40828 3596
rect 40776 3553 40785 3587
rect 40785 3553 40819 3587
rect 40819 3553 40828 3587
rect 40776 3544 40828 3553
rect 41236 3587 41288 3596
rect 41236 3553 41245 3587
rect 41245 3553 41279 3587
rect 41279 3553 41288 3587
rect 41236 3544 41288 3553
rect 46204 3587 46256 3596
rect 46204 3553 46213 3587
rect 46213 3553 46247 3587
rect 46247 3553 46256 3587
rect 46204 3544 46256 3553
rect 46388 3544 46440 3596
rect 36084 3519 36136 3528
rect 36084 3485 36093 3519
rect 36093 3485 36127 3519
rect 36127 3485 36136 3519
rect 36084 3476 36136 3485
rect 38568 3476 38620 3528
rect 29920 3340 29972 3392
rect 30288 3383 30340 3392
rect 30288 3349 30297 3383
rect 30297 3349 30331 3383
rect 30331 3349 30340 3383
rect 30288 3340 30340 3349
rect 33968 3408 34020 3460
rect 44824 3408 44876 3460
rect 47216 3408 47268 3460
rect 42524 3340 42576 3392
rect 43260 3340 43312 3392
rect 44916 3340 44968 3392
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 2136 3136 2188 3188
rect 2596 3136 2648 3188
rect 4804 3136 4856 3188
rect 2780 3068 2832 3120
rect 3700 3111 3752 3120
rect 3700 3077 3709 3111
rect 3709 3077 3743 3111
rect 3743 3077 3752 3111
rect 3700 3068 3752 3077
rect 1952 3000 2004 3052
rect 3516 3043 3568 3052
rect 3516 3009 3525 3043
rect 3525 3009 3559 3043
rect 3559 3009 3568 3043
rect 3516 3000 3568 3009
rect 2964 2932 3016 2984
rect 3240 2932 3292 2984
rect 664 2864 716 2916
rect 2688 2864 2740 2916
rect 11612 3136 11664 3188
rect 26700 3136 26752 3188
rect 30012 3136 30064 3188
rect 6276 3000 6328 3052
rect 9680 3000 9732 3052
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 11704 3000 11756 3052
rect 6644 2932 6696 2984
rect 7748 2932 7800 2984
rect 16488 3068 16540 3120
rect 17500 3111 17552 3120
rect 17500 3077 17509 3111
rect 17509 3077 17543 3111
rect 17543 3077 17552 3111
rect 17500 3068 17552 3077
rect 17684 3068 17736 3120
rect 23296 3068 23348 3120
rect 23572 3111 23624 3120
rect 23572 3077 23581 3111
rect 23581 3077 23615 3111
rect 23615 3077 23624 3111
rect 23572 3068 23624 3077
rect 25504 3068 25556 3120
rect 29460 3068 29512 3120
rect 29920 3111 29972 3120
rect 29920 3077 29926 3111
rect 29926 3077 29960 3111
rect 29960 3077 29972 3111
rect 29920 3068 29972 3077
rect 31484 3068 31536 3120
rect 34244 3136 34296 3188
rect 48044 3136 48096 3188
rect 34336 3068 34388 3120
rect 44916 3111 44968 3120
rect 15108 3000 15160 3052
rect 17316 3043 17368 3052
rect 17316 3009 17325 3043
rect 17325 3009 17359 3043
rect 17359 3009 17368 3043
rect 17316 3000 17368 3009
rect 20260 3000 20312 3052
rect 22560 3000 22612 3052
rect 23388 3043 23440 3052
rect 23388 3009 23397 3043
rect 23397 3009 23431 3043
rect 23431 3009 23440 3043
rect 23388 3000 23440 3009
rect 29552 3000 29604 3052
rect 29736 3043 29788 3052
rect 29736 3009 29745 3043
rect 29745 3009 29779 3043
rect 29779 3009 29788 3043
rect 29736 3000 29788 3009
rect 32128 3043 32180 3052
rect 32128 3009 32137 3043
rect 32137 3009 32171 3043
rect 32171 3009 32180 3043
rect 32128 3000 32180 3009
rect 36084 3000 36136 3052
rect 38568 3043 38620 3052
rect 38568 3009 38577 3043
rect 38577 3009 38611 3043
rect 38611 3009 38620 3043
rect 38568 3000 38620 3009
rect 44916 3077 44925 3111
rect 44925 3077 44959 3111
rect 44959 3077 44968 3111
rect 44916 3068 44968 3077
rect 42432 3043 42484 3052
rect 42432 3009 42441 3043
rect 42441 3009 42475 3043
rect 42475 3009 42484 3043
rect 42432 3000 42484 3009
rect 44732 3043 44784 3052
rect 44732 3009 44741 3043
rect 44741 3009 44775 3043
rect 44775 3009 44784 3043
rect 44732 3000 44784 3009
rect 49608 3000 49660 3052
rect 12440 2975 12492 2984
rect 12440 2941 12449 2975
rect 12449 2941 12483 2975
rect 12483 2941 12492 2975
rect 12440 2932 12492 2941
rect 12716 2932 12768 2984
rect 12900 2975 12952 2984
rect 12900 2941 12909 2975
rect 12909 2941 12943 2975
rect 12943 2941 12952 2975
rect 12900 2932 12952 2941
rect 7104 2864 7156 2916
rect 10968 2864 11020 2916
rect 17592 2932 17644 2984
rect 18052 2975 18104 2984
rect 18052 2941 18061 2975
rect 18061 2941 18095 2975
rect 18095 2941 18104 2975
rect 18052 2932 18104 2941
rect 23848 2975 23900 2984
rect 23848 2941 23857 2975
rect 23857 2941 23891 2975
rect 23891 2941 23900 2975
rect 23848 2932 23900 2941
rect 24124 2932 24176 2984
rect 20444 2864 20496 2916
rect 26700 2932 26752 2984
rect 31208 2932 31260 2984
rect 31300 2975 31352 2984
rect 31300 2941 31309 2975
rect 31309 2941 31343 2975
rect 31343 2941 31352 2975
rect 33508 2975 33560 2984
rect 31300 2932 31352 2941
rect 33508 2941 33517 2975
rect 33517 2941 33551 2975
rect 33551 2941 33560 2975
rect 33508 2932 33560 2941
rect 34520 2932 34572 2984
rect 38016 2932 38068 2984
rect 38752 2975 38804 2984
rect 38752 2941 38761 2975
rect 38761 2941 38795 2975
rect 38795 2941 38804 2975
rect 38752 2932 38804 2941
rect 39948 2975 40000 2984
rect 39948 2941 39957 2975
rect 39957 2941 39991 2975
rect 39991 2941 40000 2975
rect 39948 2932 40000 2941
rect 42708 2932 42760 2984
rect 45100 2932 45152 2984
rect 5816 2796 5868 2848
rect 7012 2796 7064 2848
rect 11520 2796 11572 2848
rect 18144 2796 18196 2848
rect 22744 2796 22796 2848
rect 26148 2839 26200 2848
rect 26148 2805 26157 2839
rect 26157 2805 26191 2839
rect 26191 2805 26200 2839
rect 26148 2796 26200 2805
rect 32220 2864 32272 2916
rect 41880 2796 41932 2848
rect 42708 2796 42760 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 3976 2635 4028 2644
rect 3976 2601 3985 2635
rect 3985 2601 4019 2635
rect 4019 2601 4028 2635
rect 3976 2592 4028 2601
rect 4068 2592 4120 2644
rect 9128 2592 9180 2644
rect 12440 2592 12492 2644
rect 13176 2592 13228 2644
rect 21640 2592 21692 2644
rect 46848 2592 46900 2644
rect 1308 2524 1360 2576
rect 1584 2456 1636 2508
rect 7196 2524 7248 2576
rect 20168 2524 20220 2576
rect 20352 2567 20404 2576
rect 20352 2533 20361 2567
rect 20361 2533 20395 2567
rect 20395 2533 20404 2567
rect 20352 2524 20404 2533
rect 21272 2524 21324 2576
rect 6920 2456 6972 2508
rect 7012 2499 7064 2508
rect 7012 2465 7021 2499
rect 7021 2465 7055 2499
rect 7055 2465 7064 2499
rect 7012 2456 7064 2465
rect 7472 2456 7524 2508
rect 15200 2456 15252 2508
rect 20996 2456 21048 2508
rect 24124 2524 24176 2576
rect 25872 2567 25924 2576
rect 23940 2456 23992 2508
rect 25872 2533 25881 2567
rect 25881 2533 25915 2567
rect 25915 2533 25924 2567
rect 25872 2524 25924 2533
rect 27252 2567 27304 2576
rect 27252 2533 27261 2567
rect 27261 2533 27295 2567
rect 27295 2533 27304 2567
rect 27252 2524 27304 2533
rect 30472 2524 30524 2576
rect 33140 2567 33192 2576
rect 33140 2533 33149 2567
rect 33149 2533 33183 2567
rect 33183 2533 33192 2567
rect 33140 2524 33192 2533
rect 35072 2567 35124 2576
rect 35072 2533 35081 2567
rect 35081 2533 35115 2567
rect 35115 2533 35124 2567
rect 35072 2524 35124 2533
rect 35348 2524 35400 2576
rect 38660 2524 38712 2576
rect 30288 2456 30340 2508
rect 30932 2499 30984 2508
rect 30932 2465 30941 2499
rect 30941 2465 30975 2499
rect 30975 2465 30984 2499
rect 30932 2456 30984 2465
rect 45836 2456 45888 2508
rect 4528 2388 4580 2440
rect 20536 2388 20588 2440
rect 24492 2388 24544 2440
rect 25136 2388 25188 2440
rect 27068 2431 27120 2440
rect 27068 2397 27077 2431
rect 27077 2397 27111 2431
rect 27111 2397 27120 2431
rect 27068 2388 27120 2397
rect 27712 2388 27764 2440
rect 32864 2388 32916 2440
rect 2872 2320 2924 2372
rect 8392 2320 8444 2372
rect 14188 2320 14240 2372
rect 17408 2320 17460 2372
rect 19984 2320 20036 2372
rect 21088 2320 21140 2372
rect 25780 2320 25832 2372
rect 34152 2320 34204 2372
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 10600 2295 10652 2304
rect 10600 2261 10609 2295
rect 10609 2261 10643 2295
rect 10643 2261 10652 2295
rect 10600 2252 10652 2261
rect 23020 2252 23072 2304
rect 34796 2388 34848 2440
rect 36084 2388 36136 2440
rect 38660 2388 38712 2440
rect 38108 2320 38160 2372
rect 48320 2388 48372 2440
rect 43168 2320 43220 2372
rect 46940 2320 46992 2372
rect 47768 2363 47820 2372
rect 47768 2329 47777 2363
rect 47777 2329 47811 2363
rect 47811 2329 47820 2363
rect 47768 2320 47820 2329
rect 45744 2252 45796 2304
rect 47860 2295 47912 2304
rect 47860 2261 47869 2295
rect 47869 2261 47903 2295
rect 47903 2261 47912 2295
rect 47860 2252 47912 2261
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 21824 2048 21876 2100
rect 27252 2048 27304 2100
rect 21180 1980 21232 2032
rect 33140 1980 33192 2032
rect 10600 1912 10652 1964
rect 28724 1912 28776 1964
rect 26516 1844 26568 1896
rect 47860 1844 47912 1896
rect 12256 1232 12308 1284
rect 12808 1232 12860 1284
<< metal2 >>
rect 18 51200 74 52000
rect 662 51200 718 52000
rect 1306 51200 1362 52000
rect 1950 51200 2006 52000
rect 2594 51200 2650 52000
rect 2870 51776 2926 51785
rect 2870 51711 2926 51720
rect 32 48278 60 51200
rect 676 49230 704 51200
rect 664 49224 716 49230
rect 664 49166 716 49172
rect 20 48272 72 48278
rect 20 48214 72 48220
rect 1320 48210 1348 51200
rect 1492 49088 1544 49094
rect 1492 49030 1544 49036
rect 1308 48204 1360 48210
rect 1308 48146 1360 48152
rect 1400 45960 1452 45966
rect 1400 45902 1452 45908
rect 1412 45665 1440 45902
rect 1398 45656 1454 45665
rect 1398 45591 1454 45600
rect 1400 42016 1452 42022
rect 1400 41958 1452 41964
rect 1412 41682 1440 41958
rect 1400 41676 1452 41682
rect 1400 41618 1452 41624
rect 1400 40520 1452 40526
rect 1400 40462 1452 40468
rect 1412 40225 1440 40462
rect 1398 40216 1454 40225
rect 1398 40151 1454 40160
rect 1400 37324 1452 37330
rect 1400 37266 1452 37272
rect 1412 36825 1440 37266
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1400 35080 1452 35086
rect 1400 35022 1452 35028
rect 1412 34785 1440 35022
rect 1398 34776 1454 34785
rect 1398 34711 1454 34720
rect 1400 34400 1452 34406
rect 1400 34342 1452 34348
rect 1412 34066 1440 34342
rect 1400 34060 1452 34066
rect 1400 34002 1452 34008
rect 1504 31754 1532 49030
rect 1964 48906 1992 51200
rect 2780 49156 2832 49162
rect 2780 49098 2832 49104
rect 1964 48878 2084 48906
rect 1584 48068 1636 48074
rect 1584 48010 1636 48016
rect 1596 47802 1624 48010
rect 1584 47796 1636 47802
rect 1584 47738 1636 47744
rect 1952 47592 2004 47598
rect 1952 47534 2004 47540
rect 1860 47116 1912 47122
rect 1860 47058 1912 47064
rect 1872 47025 1900 47058
rect 1858 47016 1914 47025
rect 1584 46980 1636 46986
rect 1858 46951 1914 46960
rect 1584 46922 1636 46928
rect 1596 46170 1624 46922
rect 1964 46578 1992 47534
rect 2056 46578 2084 48878
rect 2792 48278 2820 49098
rect 2884 48822 2912 51711
rect 3238 51354 3294 52000
rect 3238 51326 3648 51354
rect 3238 51200 3294 51326
rect 3620 49230 3648 51326
rect 3882 51200 3938 52000
rect 4526 51200 4582 52000
rect 5170 51354 5226 52000
rect 5170 51326 5488 51354
rect 5170 51200 5226 51326
rect 4066 51096 4122 51105
rect 4066 51031 4122 51040
rect 3974 50416 4030 50425
rect 3974 50351 4030 50360
rect 3608 49224 3660 49230
rect 3608 49166 3660 49172
rect 2964 49156 3016 49162
rect 2964 49098 3016 49104
rect 2872 48816 2924 48822
rect 2872 48758 2924 48764
rect 2780 48272 2832 48278
rect 2780 48214 2832 48220
rect 2872 47592 2924 47598
rect 2872 47534 2924 47540
rect 2884 46714 2912 47534
rect 2872 46708 2924 46714
rect 2872 46650 2924 46656
rect 1952 46572 2004 46578
rect 1952 46514 2004 46520
rect 2044 46572 2096 46578
rect 2044 46514 2096 46520
rect 2320 46572 2372 46578
rect 2320 46514 2372 46520
rect 1768 46368 1820 46374
rect 1768 46310 1820 46316
rect 1584 46164 1636 46170
rect 1584 46106 1636 46112
rect 1676 43648 1728 43654
rect 1676 43590 1728 43596
rect 1584 41540 1636 41546
rect 1584 41482 1636 41488
rect 1596 41274 1624 41482
rect 1584 41268 1636 41274
rect 1584 41210 1636 41216
rect 1584 40384 1636 40390
rect 1584 40326 1636 40332
rect 1596 35834 1624 40326
rect 1584 35828 1636 35834
rect 1584 35770 1636 35776
rect 1504 31726 1624 31754
rect 1492 31408 1544 31414
rect 1490 31376 1492 31385
rect 1544 31376 1546 31385
rect 1490 31311 1546 31320
rect 1596 30920 1624 31726
rect 1504 30892 1624 30920
rect 1400 30048 1452 30054
rect 1400 29990 1452 29996
rect 1412 29714 1440 29990
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1412 26450 1440 27406
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1400 24200 1452 24206
rect 1400 24142 1452 24148
rect 1412 23905 1440 24142
rect 1398 23896 1454 23905
rect 1398 23831 1454 23840
rect 1504 22710 1532 30892
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1596 26042 1624 26250
rect 1584 26036 1636 26042
rect 1584 25978 1636 25984
rect 1582 25936 1638 25945
rect 1582 25871 1584 25880
rect 1636 25871 1638 25880
rect 1584 25842 1636 25848
rect 1584 24064 1636 24070
rect 1584 24006 1636 24012
rect 1596 23866 1624 24006
rect 1584 23860 1636 23866
rect 1584 23802 1636 23808
rect 1492 22704 1544 22710
rect 1492 22646 1544 22652
rect 1688 22098 1716 43590
rect 1780 32910 1808 46310
rect 2332 45966 2360 46514
rect 2778 46336 2834 46345
rect 2778 46271 2834 46280
rect 2320 45960 2372 45966
rect 2320 45902 2372 45908
rect 2792 45422 2820 46271
rect 1952 45416 2004 45422
rect 1952 45358 2004 45364
rect 2780 45416 2832 45422
rect 2780 45358 2832 45364
rect 1964 44538 1992 45358
rect 2778 44976 2834 44985
rect 2778 44911 2780 44920
rect 2832 44911 2834 44920
rect 2780 44882 2832 44888
rect 2872 44736 2924 44742
rect 2872 44678 2924 44684
rect 1952 44532 2004 44538
rect 1952 44474 2004 44480
rect 1860 44396 1912 44402
rect 1860 44338 1912 44344
rect 2228 44396 2280 44402
rect 2228 44338 2280 44344
rect 1872 44305 1900 44338
rect 1858 44296 1914 44305
rect 1858 44231 1914 44240
rect 2136 44192 2188 44198
rect 2136 44134 2188 44140
rect 1860 43716 1912 43722
rect 1860 43658 1912 43664
rect 1872 43625 1900 43658
rect 1858 43616 1914 43625
rect 1858 43551 1914 43560
rect 1860 41676 1912 41682
rect 1860 41618 1912 41624
rect 1872 41585 1900 41618
rect 1858 41576 1914 41585
rect 1858 41511 1914 41520
rect 1860 41132 1912 41138
rect 1860 41074 1912 41080
rect 1872 40905 1900 41074
rect 1858 40896 1914 40905
rect 1858 40831 1914 40840
rect 2044 38888 2096 38894
rect 2044 38830 2096 38836
rect 2056 38554 2084 38830
rect 2044 38548 2096 38554
rect 2044 38490 2096 38496
rect 1860 37868 1912 37874
rect 1860 37810 1912 37816
rect 1872 37505 1900 37810
rect 1952 37664 2004 37670
rect 1952 37606 2004 37612
rect 1858 37496 1914 37505
rect 1964 37466 1992 37606
rect 1858 37431 1914 37440
rect 1952 37460 2004 37466
rect 1952 37402 2004 37408
rect 2148 37346 2176 44134
rect 1964 37318 2176 37346
rect 1964 35894 1992 37318
rect 2136 37188 2188 37194
rect 2136 37130 2188 37136
rect 2044 36576 2096 36582
rect 2044 36518 2096 36524
rect 1872 35866 1992 35894
rect 1768 32904 1820 32910
rect 1768 32846 1820 32852
rect 1768 32768 1820 32774
rect 1768 32710 1820 32716
rect 1780 32434 1808 32710
rect 1768 32428 1820 32434
rect 1768 32370 1820 32376
rect 1872 31754 1900 35866
rect 2056 35698 2084 36518
rect 2044 35692 2096 35698
rect 2044 35634 2096 35640
rect 2148 34082 2176 37130
rect 2056 34054 2176 34082
rect 1952 32360 2004 32366
rect 1952 32302 2004 32308
rect 1780 31726 1900 31754
rect 1780 27554 1808 31726
rect 1964 30938 1992 32302
rect 2056 31754 2084 34054
rect 2136 33924 2188 33930
rect 2136 33866 2188 33872
rect 2148 33658 2176 33866
rect 2136 33652 2188 33658
rect 2136 33594 2188 33600
rect 2240 33522 2268 44338
rect 2884 43994 2912 44678
rect 2872 43988 2924 43994
rect 2872 43930 2924 43936
rect 2976 41138 3004 49098
rect 3146 49056 3202 49065
rect 3146 48991 3202 49000
rect 3056 48680 3108 48686
rect 3056 48622 3108 48628
rect 3068 47258 3096 48622
rect 3160 47598 3188 48991
rect 3422 48376 3478 48385
rect 3422 48311 3424 48320
rect 3476 48311 3478 48320
rect 3424 48282 3476 48288
rect 3988 48278 4016 50351
rect 4080 49774 4108 51031
rect 4068 49768 4120 49774
rect 4068 49710 4120 49716
rect 4540 49722 4568 51200
rect 4540 49694 4660 49722
rect 4214 49532 4522 49552
rect 4214 49530 4220 49532
rect 4276 49530 4300 49532
rect 4356 49530 4380 49532
rect 4436 49530 4460 49532
rect 4516 49530 4522 49532
rect 4276 49478 4278 49530
rect 4458 49478 4460 49530
rect 4214 49476 4220 49478
rect 4276 49476 4300 49478
rect 4356 49476 4380 49478
rect 4436 49476 4460 49478
rect 4516 49476 4522 49478
rect 4214 49456 4522 49476
rect 4632 49230 4660 49694
rect 4620 49224 4672 49230
rect 4620 49166 4672 49172
rect 4620 49088 4672 49094
rect 4620 49030 4672 49036
rect 5264 49088 5316 49094
rect 5264 49030 5316 49036
rect 4214 48444 4522 48464
rect 4214 48442 4220 48444
rect 4276 48442 4300 48444
rect 4356 48442 4380 48444
rect 4436 48442 4460 48444
rect 4516 48442 4522 48444
rect 4276 48390 4278 48442
rect 4458 48390 4460 48442
rect 4214 48388 4220 48390
rect 4276 48388 4300 48390
rect 4356 48388 4380 48390
rect 4436 48388 4460 48390
rect 4516 48388 4522 48390
rect 4214 48368 4522 48388
rect 3976 48272 4028 48278
rect 3976 48214 4028 48220
rect 3792 48136 3844 48142
rect 3792 48078 3844 48084
rect 3804 47705 3832 48078
rect 3884 48000 3936 48006
rect 3884 47942 3936 47948
rect 4068 48000 4120 48006
rect 4068 47942 4120 47948
rect 3790 47696 3846 47705
rect 3790 47631 3846 47640
rect 3148 47592 3200 47598
rect 3148 47534 3200 47540
rect 3056 47252 3108 47258
rect 3056 47194 3108 47200
rect 3608 47184 3660 47190
rect 3608 47126 3660 47132
rect 3332 47048 3384 47054
rect 3332 46990 3384 46996
rect 3148 45960 3200 45966
rect 3148 45902 3200 45908
rect 3160 45558 3188 45902
rect 3148 45552 3200 45558
rect 3148 45494 3200 45500
rect 3344 44402 3372 46990
rect 3620 46578 3648 47126
rect 3608 46572 3660 46578
rect 3608 46514 3660 46520
rect 3896 46170 3924 47942
rect 3884 46164 3936 46170
rect 3884 46106 3936 46112
rect 3424 44804 3476 44810
rect 3424 44746 3476 44752
rect 3436 44538 3464 44746
rect 3424 44532 3476 44538
rect 3424 44474 3476 44480
rect 3332 44396 3384 44402
rect 3332 44338 3384 44344
rect 2320 41132 2372 41138
rect 2320 41074 2372 41080
rect 2964 41132 3016 41138
rect 2964 41074 3016 41080
rect 2332 37194 2360 41074
rect 2412 40996 2464 41002
rect 2412 40938 2464 40944
rect 2320 37188 2372 37194
rect 2320 37130 2372 37136
rect 2424 35894 2452 40938
rect 2870 39536 2926 39545
rect 2870 39471 2926 39480
rect 2884 38894 2912 39471
rect 2780 38888 2832 38894
rect 2780 38830 2832 38836
rect 2872 38888 2924 38894
rect 2872 38830 2924 38836
rect 2792 38010 2820 38830
rect 2780 38004 2832 38010
rect 2780 37946 2832 37952
rect 3344 36378 3372 44338
rect 4080 41414 4108 47942
rect 4214 47356 4522 47376
rect 4214 47354 4220 47356
rect 4276 47354 4300 47356
rect 4356 47354 4380 47356
rect 4436 47354 4460 47356
rect 4516 47354 4522 47356
rect 4276 47302 4278 47354
rect 4458 47302 4460 47354
rect 4214 47300 4220 47302
rect 4276 47300 4300 47302
rect 4356 47300 4380 47302
rect 4436 47300 4460 47302
rect 4516 47300 4522 47302
rect 4214 47280 4522 47300
rect 4214 46268 4522 46288
rect 4214 46266 4220 46268
rect 4276 46266 4300 46268
rect 4356 46266 4380 46268
rect 4436 46266 4460 46268
rect 4516 46266 4522 46268
rect 4276 46214 4278 46266
rect 4458 46214 4460 46266
rect 4214 46212 4220 46214
rect 4276 46212 4300 46214
rect 4356 46212 4380 46214
rect 4436 46212 4460 46214
rect 4516 46212 4522 46214
rect 4214 46192 4522 46212
rect 4214 45180 4522 45200
rect 4214 45178 4220 45180
rect 4276 45178 4300 45180
rect 4356 45178 4380 45180
rect 4436 45178 4460 45180
rect 4516 45178 4522 45180
rect 4276 45126 4278 45178
rect 4458 45126 4460 45178
rect 4214 45124 4220 45126
rect 4276 45124 4300 45126
rect 4356 45124 4380 45126
rect 4436 45124 4460 45126
rect 4516 45124 4522 45126
rect 4214 45104 4522 45124
rect 4214 44092 4522 44112
rect 4214 44090 4220 44092
rect 4276 44090 4300 44092
rect 4356 44090 4380 44092
rect 4436 44090 4460 44092
rect 4516 44090 4522 44092
rect 4276 44038 4278 44090
rect 4458 44038 4460 44090
rect 4214 44036 4220 44038
rect 4276 44036 4300 44038
rect 4356 44036 4380 44038
rect 4436 44036 4460 44038
rect 4516 44036 4522 44038
rect 4214 44016 4522 44036
rect 4214 43004 4522 43024
rect 4214 43002 4220 43004
rect 4276 43002 4300 43004
rect 4356 43002 4380 43004
rect 4436 43002 4460 43004
rect 4516 43002 4522 43004
rect 4276 42950 4278 43002
rect 4458 42950 4460 43002
rect 4214 42948 4220 42950
rect 4276 42948 4300 42950
rect 4356 42948 4380 42950
rect 4436 42948 4460 42950
rect 4516 42948 4522 42950
rect 4214 42928 4522 42948
rect 4214 41916 4522 41936
rect 4214 41914 4220 41916
rect 4276 41914 4300 41916
rect 4356 41914 4380 41916
rect 4436 41914 4460 41916
rect 4516 41914 4522 41916
rect 4276 41862 4278 41914
rect 4458 41862 4460 41914
rect 4214 41860 4220 41862
rect 4276 41860 4300 41862
rect 4356 41860 4380 41862
rect 4436 41860 4460 41862
rect 4516 41860 4522 41862
rect 4214 41840 4522 41860
rect 3988 41386 4108 41414
rect 3988 37210 4016 41386
rect 4214 40828 4522 40848
rect 4214 40826 4220 40828
rect 4276 40826 4300 40828
rect 4356 40826 4380 40828
rect 4436 40826 4460 40828
rect 4516 40826 4522 40828
rect 4276 40774 4278 40826
rect 4458 40774 4460 40826
rect 4214 40772 4220 40774
rect 4276 40772 4300 40774
rect 4356 40772 4380 40774
rect 4436 40772 4460 40774
rect 4516 40772 4522 40774
rect 4214 40752 4522 40772
rect 4214 39740 4522 39760
rect 4214 39738 4220 39740
rect 4276 39738 4300 39740
rect 4356 39738 4380 39740
rect 4436 39738 4460 39740
rect 4516 39738 4522 39740
rect 4276 39686 4278 39738
rect 4458 39686 4460 39738
rect 4214 39684 4220 39686
rect 4276 39684 4300 39686
rect 4356 39684 4380 39686
rect 4436 39684 4460 39686
rect 4516 39684 4522 39686
rect 4214 39664 4522 39684
rect 4214 38652 4522 38672
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38576 4522 38596
rect 4066 38176 4122 38185
rect 4066 38111 4122 38120
rect 4080 37330 4108 38111
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 4068 37324 4120 37330
rect 4068 37266 4120 37272
rect 3988 37182 4108 37210
rect 3332 36372 3384 36378
rect 3332 36314 3384 36320
rect 3332 36168 3384 36174
rect 2778 36136 2834 36145
rect 3332 36110 3384 36116
rect 2778 36071 2834 36080
rect 2424 35866 2544 35894
rect 2228 33516 2280 33522
rect 2228 33458 2280 33464
rect 2056 31726 2176 31754
rect 1952 30932 2004 30938
rect 1952 30874 2004 30880
rect 2044 30252 2096 30258
rect 2044 30194 2096 30200
rect 1860 28960 1912 28966
rect 1860 28902 1912 28908
rect 1872 28626 1900 28902
rect 1860 28620 1912 28626
rect 1860 28562 1912 28568
rect 1780 27526 1900 27554
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1780 26994 1808 27338
rect 1768 26988 1820 26994
rect 1768 26930 1820 26936
rect 1872 26874 1900 27526
rect 1952 27328 2004 27334
rect 1952 27270 2004 27276
rect 1964 27062 1992 27270
rect 1952 27056 2004 27062
rect 1952 26998 2004 27004
rect 1780 26846 1900 26874
rect 1676 22092 1728 22098
rect 1676 22034 1728 22040
rect 1584 18080 1636 18086
rect 1584 18022 1636 18028
rect 1596 17746 1624 18022
rect 1584 17740 1636 17746
rect 1584 17682 1636 17688
rect 1400 17128 1452 17134
rect 1400 17070 1452 17076
rect 1412 16794 1440 17070
rect 1780 16998 1808 26846
rect 2056 25158 2084 30194
rect 2044 25152 2096 25158
rect 2044 25094 2096 25100
rect 2056 24426 2084 25094
rect 1964 24398 2084 24426
rect 1860 22636 1912 22642
rect 1860 22578 1912 22584
rect 1872 22545 1900 22578
rect 1964 22574 1992 24398
rect 2044 23520 2096 23526
rect 2044 23462 2096 23468
rect 2056 23186 2084 23462
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 1952 22568 2004 22574
rect 1858 22536 1914 22545
rect 1952 22510 2004 22516
rect 1858 22471 1914 22480
rect 1952 22432 2004 22438
rect 1952 22374 2004 22380
rect 1964 22234 1992 22374
rect 1952 22228 2004 22234
rect 1952 22170 2004 22176
rect 1860 19848 1912 19854
rect 1860 19790 1912 19796
rect 1872 19378 1900 19790
rect 1860 19372 1912 19378
rect 1860 19314 1912 19320
rect 2044 19304 2096 19310
rect 2044 19246 2096 19252
rect 2056 18970 2084 19246
rect 2044 18964 2096 18970
rect 2044 18906 2096 18912
rect 2148 18850 2176 31726
rect 2240 27470 2268 33458
rect 2320 30048 2372 30054
rect 2320 29990 2372 29996
rect 2332 29714 2360 29990
rect 2320 29708 2372 29714
rect 2320 29650 2372 29656
rect 2412 28960 2464 28966
rect 2412 28902 2464 28908
rect 2424 28490 2452 28902
rect 2412 28484 2464 28490
rect 2412 28426 2464 28432
rect 2516 27690 2544 35866
rect 2792 35630 2820 36071
rect 3056 36032 3108 36038
rect 3056 35974 3108 35980
rect 3068 35766 3096 35974
rect 3056 35760 3108 35766
rect 3056 35702 3108 35708
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2778 34096 2834 34105
rect 2778 34031 2780 34040
rect 2832 34031 2834 34040
rect 2780 34002 2832 34008
rect 2778 33416 2834 33425
rect 2778 33351 2834 33360
rect 2596 32904 2648 32910
rect 2596 32846 2648 32852
rect 2332 27662 2544 27690
rect 2228 27464 2280 27470
rect 2228 27406 2280 27412
rect 2240 26246 2268 27406
rect 2228 26240 2280 26246
rect 2228 26182 2280 26188
rect 2228 25900 2280 25906
rect 2228 25842 2280 25848
rect 2240 24614 2268 25842
rect 2228 24608 2280 24614
rect 2228 24550 2280 24556
rect 2056 18822 2176 18850
rect 1858 17096 1914 17105
rect 1858 17031 1914 17040
rect 1768 16992 1820 16998
rect 1768 16934 1820 16940
rect 1400 16788 1452 16794
rect 1400 16730 1452 16736
rect 1872 16590 1900 17031
rect 1860 16584 1912 16590
rect 2056 16574 2084 18822
rect 2136 18080 2188 18086
rect 2136 18022 2188 18028
rect 2148 17610 2176 18022
rect 2136 17604 2188 17610
rect 2136 17546 2188 17552
rect 2056 16546 2176 16574
rect 1860 16526 1912 16532
rect 20 16448 72 16454
rect 20 16390 72 16396
rect 32 800 60 16390
rect 1768 14408 1820 14414
rect 1768 14350 1820 14356
rect 1780 13938 1808 14350
rect 1768 13932 1820 13938
rect 1768 13874 1820 13880
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13530 1992 13806
rect 1952 13524 2004 13530
rect 1952 13466 2004 13472
rect 1952 13320 2004 13326
rect 1952 13262 2004 13268
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 12345 1440 12718
rect 1398 12336 1454 12345
rect 1398 12271 1454 12280
rect 1584 11552 1636 11558
rect 1584 11494 1636 11500
rect 1398 10976 1454 10985
rect 1398 10911 1454 10920
rect 1412 10674 1440 10911
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1596 9994 1624 11494
rect 1584 9988 1636 9994
rect 1584 9930 1636 9936
rect 1860 8492 1912 8498
rect 1860 8434 1912 8440
rect 1872 8265 1900 8434
rect 1858 8256 1914 8265
rect 1858 8191 1914 8200
rect 1860 7812 1912 7818
rect 1860 7754 1912 7760
rect 1872 7585 1900 7754
rect 1858 7576 1914 7585
rect 1858 7511 1914 7520
rect 1400 5024 1452 5030
rect 1400 4966 1452 4972
rect 1412 4690 1440 4966
rect 1400 4684 1452 4690
rect 1400 4626 1452 4632
rect 1964 4146 1992 13262
rect 2044 7200 2096 7206
rect 2044 7142 2096 7148
rect 2056 6866 2084 7142
rect 2044 6860 2096 6866
rect 2044 6802 2096 6808
rect 2148 6322 2176 16546
rect 2240 11762 2268 24550
rect 2332 23594 2360 27662
rect 2608 26908 2636 32846
rect 2792 32366 2820 33351
rect 2872 33312 2924 33318
rect 2872 33254 2924 33260
rect 2780 32360 2832 32366
rect 2780 32302 2832 32308
rect 2884 31210 2912 33254
rect 3056 32768 3108 32774
rect 3056 32710 3108 32716
rect 3146 32736 3202 32745
rect 2964 31952 3016 31958
rect 2964 31894 3016 31900
rect 2872 31204 2924 31210
rect 2872 31146 2924 31152
rect 2976 30938 3004 31894
rect 3068 31414 3096 32710
rect 3146 32671 3202 32680
rect 3056 31408 3108 31414
rect 3056 31350 3108 31356
rect 3160 31278 3188 32671
rect 3238 32056 3294 32065
rect 3238 31991 3294 32000
rect 3252 31822 3280 31991
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 3148 31272 3200 31278
rect 3148 31214 3200 31220
rect 2964 30932 3016 30938
rect 2964 30874 3016 30880
rect 2964 30728 3016 30734
rect 2964 30670 3016 30676
rect 2778 30016 2834 30025
rect 2778 29951 2834 29960
rect 2792 29714 2820 29951
rect 2780 29708 2832 29714
rect 2780 29650 2832 29656
rect 2976 29170 3004 30670
rect 2688 29164 2740 29170
rect 2688 29106 2740 29112
rect 2964 29164 3016 29170
rect 2964 29106 3016 29112
rect 2424 26880 2636 26908
rect 2320 23588 2372 23594
rect 2320 23530 2372 23536
rect 2424 21554 2452 26880
rect 2700 23526 2728 29106
rect 2872 28960 2924 28966
rect 2872 28902 2924 28908
rect 2778 28656 2834 28665
rect 2778 28591 2780 28600
rect 2832 28591 2834 28600
rect 2780 28562 2832 28568
rect 2884 28150 2912 28902
rect 2872 28144 2924 28150
rect 2872 28086 2924 28092
rect 2778 27296 2834 27305
rect 2778 27231 2834 27240
rect 2792 26926 2820 27231
rect 2780 26920 2832 26926
rect 2780 26862 2832 26868
rect 2778 26616 2834 26625
rect 2778 26551 2834 26560
rect 2792 26450 2820 26551
rect 2780 26444 2832 26450
rect 2780 26386 2832 26392
rect 2976 26042 3004 29106
rect 3344 27402 3372 36110
rect 3976 32904 4028 32910
rect 3976 32846 4028 32852
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3332 27396 3384 27402
rect 3332 27338 3384 27344
rect 3804 26586 3832 31758
rect 3792 26580 3844 26586
rect 3792 26522 3844 26528
rect 3988 26314 4016 32846
rect 4080 32026 4108 37182
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4068 32020 4120 32026
rect 4068 31962 4120 31968
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4066 29336 4122 29345
rect 4066 29271 4122 29280
rect 4080 28642 4108 29271
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4080 28614 4200 28642
rect 4172 28014 4200 28614
rect 4160 28008 4212 28014
rect 4160 27950 4212 27956
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 3976 26308 4028 26314
rect 3976 26250 4028 26256
rect 2964 26036 3016 26042
rect 2964 25978 3016 25984
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 2688 23520 2740 23526
rect 2688 23462 2740 23468
rect 2504 23248 2556 23254
rect 2504 23190 2556 23196
rect 2516 22642 2544 23190
rect 2596 23044 2648 23050
rect 2596 22986 2648 22992
rect 2608 22778 2636 22986
rect 2596 22772 2648 22778
rect 2596 22714 2648 22720
rect 2504 22636 2556 22642
rect 2504 22578 2556 22584
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2332 13326 2360 18158
rect 2320 13320 2372 13326
rect 2320 13262 2372 13268
rect 2228 11756 2280 11762
rect 2228 11698 2280 11704
rect 2228 6724 2280 6730
rect 2228 6666 2280 6672
rect 2240 6458 2268 6666
rect 2228 6452 2280 6458
rect 2228 6394 2280 6400
rect 2136 6316 2188 6322
rect 2136 6258 2188 6264
rect 2136 5704 2188 5710
rect 2136 5646 2188 5652
rect 2148 5234 2176 5646
rect 2136 5228 2188 5234
rect 2136 5170 2188 5176
rect 1952 4140 2004 4146
rect 1952 4082 2004 4088
rect 2136 4072 2188 4078
rect 2136 4014 2188 4020
rect 1584 3936 1636 3942
rect 1584 3878 1636 3884
rect 1676 3936 1728 3942
rect 1676 3878 1728 3884
rect 664 2916 716 2922
rect 664 2858 716 2864
rect 676 800 704 2858
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1320 800 1348 2518
rect 1596 2514 1624 3878
rect 1688 3602 1716 3878
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 1860 3596 1912 3602
rect 1860 3538 1912 3544
rect 1872 3505 1900 3538
rect 1858 3496 1914 3505
rect 1858 3431 1914 3440
rect 2148 3194 2176 4014
rect 2516 4010 2544 22578
rect 2596 22568 2648 22574
rect 2596 22510 2648 22516
rect 2608 16574 2636 22510
rect 2700 18290 2728 23462
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 2778 23216 2834 23225
rect 2778 23151 2780 23160
rect 2832 23151 2834 23160
rect 2780 23122 2832 23128
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3974 21856 4030 21865
rect 3974 21791 4030 21800
rect 3988 21078 4016 21791
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4066 21176 4122 21185
rect 4214 21168 4522 21188
rect 4632 21146 4660 49030
rect 4896 48680 4948 48686
rect 4896 48622 4948 48628
rect 4712 48612 4764 48618
rect 4712 48554 4764 48560
rect 4724 46578 4752 48554
rect 4804 47660 4856 47666
rect 4804 47602 4856 47608
rect 4712 46572 4764 46578
rect 4712 46514 4764 46520
rect 4816 45554 4844 47602
rect 4908 47258 4936 48622
rect 4988 48068 5040 48074
rect 4988 48010 5040 48016
rect 5000 47802 5028 48010
rect 4988 47796 5040 47802
rect 4988 47738 5040 47744
rect 4896 47252 4948 47258
rect 4896 47194 4948 47200
rect 4724 45526 4844 45554
rect 4724 23254 4752 45526
rect 5276 31414 5304 49030
rect 5460 48906 5488 51326
rect 5814 51200 5870 52000
rect 6458 51354 6514 52000
rect 6196 51326 6514 51354
rect 5632 49768 5684 49774
rect 5632 49710 5684 49716
rect 5460 48878 5580 48906
rect 5552 48822 5580 48878
rect 5540 48816 5592 48822
rect 5540 48758 5592 48764
rect 5644 48686 5672 49710
rect 5632 48680 5684 48686
rect 5632 48622 5684 48628
rect 5356 48544 5408 48550
rect 5356 48486 5408 48492
rect 5368 46578 5396 48486
rect 5540 48204 5592 48210
rect 5540 48146 5592 48152
rect 5552 47258 5580 48146
rect 6196 47734 6224 51326
rect 6458 51200 6514 51326
rect 7102 51200 7158 52000
rect 7746 51200 7802 52000
rect 8390 51354 8446 52000
rect 8312 51326 8446 51354
rect 7116 49298 7144 51200
rect 7760 49298 7788 51200
rect 6920 49292 6972 49298
rect 6920 49234 6972 49240
rect 7104 49292 7156 49298
rect 7104 49234 7156 49240
rect 7748 49292 7800 49298
rect 7748 49234 7800 49240
rect 6368 48680 6420 48686
rect 6368 48622 6420 48628
rect 6184 47728 6236 47734
rect 6184 47670 6236 47676
rect 6092 47660 6144 47666
rect 6092 47602 6144 47608
rect 5540 47252 5592 47258
rect 5540 47194 5592 47200
rect 6104 47054 6132 47602
rect 6092 47048 6144 47054
rect 6092 46990 6144 46996
rect 5356 46572 5408 46578
rect 5356 46514 5408 46520
rect 5264 31408 5316 31414
rect 5264 31350 5316 31356
rect 6380 29782 6408 48622
rect 6644 48340 6696 48346
rect 6644 48282 6696 48288
rect 6656 47598 6684 48282
rect 6552 47592 6604 47598
rect 6552 47534 6604 47540
rect 6644 47592 6696 47598
rect 6644 47534 6696 47540
rect 6564 47258 6592 47534
rect 6644 47456 6696 47462
rect 6644 47398 6696 47404
rect 6552 47252 6604 47258
rect 6552 47194 6604 47200
rect 6368 29776 6420 29782
rect 6368 29718 6420 29724
rect 6552 27056 6604 27062
rect 6552 26998 6604 27004
rect 4804 26512 4856 26518
rect 4804 26454 4856 26460
rect 4712 23248 4764 23254
rect 4712 23190 4764 23196
rect 4066 21111 4122 21120
rect 4620 21140 4672 21146
rect 3976 21072 4028 21078
rect 3976 21014 4028 21020
rect 4080 21010 4108 21111
rect 4620 21082 4672 21088
rect 4068 21004 4120 21010
rect 4068 20946 4120 20952
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 4080 19718 4108 19751
rect 4068 19712 4120 19718
rect 4068 19654 4120 19660
rect 2780 19304 2832 19310
rect 2780 19246 2832 19252
rect 2792 19145 2820 19246
rect 3516 19236 3568 19242
rect 3516 19178 3568 19184
rect 2778 19136 2834 19145
rect 2778 19071 2834 19080
rect 3146 18456 3202 18465
rect 3146 18391 3202 18400
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 3160 18154 3188 18391
rect 3148 18148 3200 18154
rect 3148 18090 3200 18096
rect 2872 18080 2924 18086
rect 2872 18022 2924 18028
rect 2778 17776 2834 17785
rect 2778 17711 2780 17720
rect 2832 17711 2834 17720
rect 2780 17682 2832 17688
rect 2884 17270 2912 18022
rect 2872 17264 2924 17270
rect 2872 17206 2924 17212
rect 2780 17128 2832 17134
rect 2780 17070 2832 17076
rect 2608 16546 2728 16574
rect 2700 4146 2728 16546
rect 2792 16425 2820 17070
rect 2778 16416 2834 16425
rect 2778 16351 2834 16360
rect 2780 13864 2832 13870
rect 2780 13806 2832 13812
rect 2792 13705 2820 13806
rect 2778 13696 2834 13705
rect 2778 13631 2834 13640
rect 3528 12850 3556 19178
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 3792 18828 3844 18834
rect 3792 18770 3844 18776
rect 3516 12844 3568 12850
rect 3516 12786 3568 12792
rect 2964 11552 3016 11558
rect 2964 11494 3016 11500
rect 2976 11218 3004 11494
rect 2964 11212 3016 11218
rect 2964 11154 3016 11160
rect 3056 11212 3108 11218
rect 3056 11154 3108 11160
rect 2872 11076 2924 11082
rect 2872 11018 2924 11024
rect 2884 10606 2912 11018
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 3068 10305 3096 11154
rect 3516 10464 3568 10470
rect 3516 10406 3568 10412
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 3528 10130 3556 10406
rect 3516 10124 3568 10130
rect 3516 10066 3568 10072
rect 3240 9988 3292 9994
rect 3240 9930 3292 9936
rect 2964 9648 3016 9654
rect 3252 9625 3280 9930
rect 2964 9590 3016 9596
rect 3238 9616 3294 9625
rect 2976 8945 3004 9590
rect 3238 9551 3294 9560
rect 2962 8936 3018 8945
rect 2962 8871 3018 8880
rect 2778 6896 2834 6905
rect 2778 6831 2780 6840
rect 2832 6831 2834 6840
rect 2780 6802 2832 6808
rect 3422 6216 3478 6225
rect 3422 6151 3478 6160
rect 3436 5914 3464 6151
rect 3424 5908 3476 5914
rect 3424 5850 3476 5856
rect 3056 5568 3108 5574
rect 2778 5536 2834 5545
rect 3056 5510 3108 5516
rect 2778 5471 2834 5480
rect 2792 5166 2820 5471
rect 3068 5302 3096 5510
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 2780 5160 2832 5166
rect 2780 5102 2832 5108
rect 3238 4856 3294 4865
rect 3238 4791 3294 4800
rect 3252 4622 3280 4791
rect 3804 4622 3832 18770
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 3884 17128 3936 17134
rect 3884 17070 3936 17076
rect 4068 17128 4120 17134
rect 4068 17070 4120 17076
rect 3896 16794 3924 17070
rect 3884 16788 3936 16794
rect 3884 16730 3936 16736
rect 4080 13025 4108 17070
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4066 13016 4122 13025
rect 4066 12951 4122 12960
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3240 4616 3292 4622
rect 3240 4558 3292 4564
rect 3792 4616 3844 4622
rect 3792 4558 3844 4564
rect 3424 4208 3476 4214
rect 3422 4176 3424 4185
rect 3476 4176 3478 4185
rect 2688 4140 2740 4146
rect 3422 4111 3478 4120
rect 2688 4082 2740 4088
rect 2504 4004 2556 4010
rect 2504 3946 2556 3952
rect 2136 3188 2188 3194
rect 2136 3130 2188 3136
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 1584 2508 1636 2514
rect 1584 2450 1636 2456
rect 1964 800 1992 2994
rect 2608 800 2636 3130
rect 2700 2922 2728 4082
rect 2872 3936 2924 3942
rect 2872 3878 2924 3884
rect 3516 3936 3568 3942
rect 3516 3878 3568 3884
rect 2780 3120 2832 3126
rect 2780 3062 2832 3068
rect 2688 2916 2740 2922
rect 2688 2858 2740 2864
rect 18 0 74 800
rect 662 0 718 800
rect 1306 0 1362 800
rect 1950 0 2006 800
rect 2594 0 2650 800
rect 2792 785 2820 3062
rect 2884 2378 2912 3878
rect 2964 3732 3016 3738
rect 2964 3674 3016 3680
rect 2976 2990 3004 3674
rect 3528 3058 3556 3878
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 3884 3528 3936 3534
rect 3884 3470 3936 3476
rect 3700 3392 3752 3398
rect 3700 3334 3752 3340
rect 3712 3126 3740 3334
rect 3700 3120 3752 3126
rect 3700 3062 3752 3068
rect 3516 3052 3568 3058
rect 3516 2994 3568 3000
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 3240 2984 3292 2990
rect 3240 2926 3292 2932
rect 2872 2372 2924 2378
rect 2872 2314 2924 2320
rect 3252 800 3280 2926
rect 3896 800 3924 3470
rect 3976 3460 4028 3466
rect 3976 3402 4028 3408
rect 3988 2650 4016 3402
rect 4816 3194 4844 26454
rect 6564 26450 6592 26998
rect 6552 26444 6604 26450
rect 6552 26386 6604 26392
rect 6656 25906 6684 47398
rect 6932 47258 6960 49234
rect 7380 49156 7432 49162
rect 7380 49098 7432 49104
rect 7392 48278 7420 49098
rect 7564 48680 7616 48686
rect 7564 48622 7616 48628
rect 7576 48278 7604 48622
rect 7380 48272 7432 48278
rect 7380 48214 7432 48220
rect 7564 48272 7616 48278
rect 7564 48214 7616 48220
rect 7196 48136 7248 48142
rect 7196 48078 7248 48084
rect 7932 48136 7984 48142
rect 7932 48078 7984 48084
rect 6920 47252 6972 47258
rect 6920 47194 6972 47200
rect 6920 28076 6972 28082
rect 6920 28018 6972 28024
rect 6932 27470 6960 28018
rect 7012 27940 7064 27946
rect 7012 27882 7064 27888
rect 6920 27464 6972 27470
rect 6920 27406 6972 27412
rect 6736 26784 6788 26790
rect 6736 26726 6788 26732
rect 6748 26450 6776 26726
rect 6736 26444 6788 26450
rect 6736 26386 6788 26392
rect 6644 25900 6696 25906
rect 6644 25842 6696 25848
rect 6276 25832 6328 25838
rect 6276 25774 6328 25780
rect 6288 6914 6316 25774
rect 6828 25696 6880 25702
rect 6828 25638 6880 25644
rect 6840 25498 6868 25638
rect 6828 25492 6880 25498
rect 6828 25434 6880 25440
rect 7024 22030 7052 27882
rect 7208 26994 7236 48078
rect 7944 47054 7972 48078
rect 7748 47048 7800 47054
rect 7748 46990 7800 46996
rect 7932 47048 7984 47054
rect 7932 46990 7984 46996
rect 7760 43790 7788 46990
rect 7748 43784 7800 43790
rect 7748 43726 7800 43732
rect 7288 37868 7340 37874
rect 7288 37810 7340 37816
rect 7300 37262 7328 37810
rect 7288 37256 7340 37262
rect 7288 37198 7340 37204
rect 7196 26988 7248 26994
rect 7196 26930 7248 26936
rect 7300 24070 7328 37198
rect 7380 37120 7432 37126
rect 7380 37062 7432 37068
rect 7392 36854 7420 37062
rect 7380 36848 7432 36854
rect 7380 36790 7432 36796
rect 7656 36100 7708 36106
rect 7656 36042 7708 36048
rect 7668 35834 7696 36042
rect 7656 35828 7708 35834
rect 7656 35770 7708 35776
rect 7380 26920 7432 26926
rect 7380 26862 7432 26868
rect 7288 24064 7340 24070
rect 7288 24006 7340 24012
rect 7392 23730 7420 26862
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7564 24812 7616 24818
rect 7564 24754 7616 24760
rect 7656 24812 7708 24818
rect 7656 24754 7708 24760
rect 7576 24342 7604 24754
rect 7564 24336 7616 24342
rect 7564 24278 7616 24284
rect 7668 24138 7696 24754
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7380 23724 7432 23730
rect 7380 23666 7432 23672
rect 7564 23656 7616 23662
rect 7564 23598 7616 23604
rect 7576 23322 7604 23598
rect 7564 23316 7616 23322
rect 7564 23258 7616 23264
rect 7760 23118 7788 25842
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7944 22094 7972 46990
rect 8312 41414 8340 51326
rect 8390 51200 8446 51326
rect 9034 51200 9090 52000
rect 9678 51200 9734 52000
rect 10322 51200 10378 52000
rect 10966 51200 11022 52000
rect 11610 51200 11666 52000
rect 12254 51354 12310 52000
rect 12898 51354 12954 52000
rect 12254 51326 12388 51354
rect 12254 51200 12310 51326
rect 8944 49224 8996 49230
rect 8944 49166 8996 49172
rect 8484 49156 8536 49162
rect 8484 49098 8536 49104
rect 8496 47258 8524 49098
rect 8956 47666 8984 49166
rect 9692 48686 9720 51200
rect 9128 48680 9180 48686
rect 9128 48622 9180 48628
rect 9680 48680 9732 48686
rect 9680 48622 9732 48628
rect 9140 48210 9168 48622
rect 9128 48204 9180 48210
rect 9128 48146 9180 48152
rect 10336 48074 10364 51200
rect 10508 48816 10560 48822
rect 10508 48758 10560 48764
rect 10048 48068 10100 48074
rect 10048 48010 10100 48016
rect 10324 48068 10376 48074
rect 10324 48010 10376 48016
rect 10060 47802 10088 48010
rect 10520 47802 10548 48758
rect 10048 47796 10100 47802
rect 10048 47738 10100 47744
rect 10508 47796 10560 47802
rect 10508 47738 10560 47744
rect 8944 47660 8996 47666
rect 8944 47602 8996 47608
rect 10980 47258 11008 51200
rect 11624 49230 11652 51200
rect 11612 49224 11664 49230
rect 11612 49166 11664 49172
rect 12072 49088 12124 49094
rect 12072 49030 12124 49036
rect 11704 48544 11756 48550
rect 11704 48486 11756 48492
rect 11716 48210 11744 48486
rect 11704 48204 11756 48210
rect 11704 48146 11756 48152
rect 8484 47252 8536 47258
rect 8484 47194 8536 47200
rect 10968 47252 11020 47258
rect 10968 47194 11020 47200
rect 11520 46640 11572 46646
rect 11520 46582 11572 46588
rect 8312 41386 8432 41414
rect 8300 37324 8352 37330
rect 8300 37266 8352 37272
rect 8312 36718 8340 37266
rect 8208 36712 8260 36718
rect 8208 36654 8260 36660
rect 8300 36712 8352 36718
rect 8300 36654 8352 36660
rect 8220 36378 8248 36654
rect 8208 36372 8260 36378
rect 8208 36314 8260 36320
rect 8404 35834 8432 41386
rect 8392 35828 8444 35834
rect 8392 35770 8444 35776
rect 11532 34610 11560 46582
rect 12084 41414 12112 49030
rect 12360 48906 12388 51326
rect 12728 51326 12954 51354
rect 12728 49298 12756 51326
rect 12898 51200 12954 51326
rect 13542 51354 13598 52000
rect 14186 51354 14242 52000
rect 14830 51354 14886 52000
rect 15474 51354 15530 52000
rect 13542 51326 13768 51354
rect 13542 51200 13598 51326
rect 13740 49314 13768 51326
rect 14186 51326 14504 51354
rect 14186 51200 14242 51326
rect 12716 49292 12768 49298
rect 13740 49286 13860 49314
rect 14476 49298 14504 51326
rect 14830 51326 15056 51354
rect 14830 51200 14886 51326
rect 12716 49234 12768 49240
rect 13832 49230 13860 49286
rect 14464 49292 14516 49298
rect 14464 49234 14516 49240
rect 13820 49224 13872 49230
rect 13820 49166 13872 49172
rect 14648 49088 14700 49094
rect 14648 49030 14700 49036
rect 12360 48878 12572 48906
rect 12440 48680 12492 48686
rect 12440 48622 12492 48628
rect 12452 48346 12480 48622
rect 12544 48618 12572 48878
rect 12808 48680 12860 48686
rect 12808 48622 12860 48628
rect 12532 48612 12584 48618
rect 12532 48554 12584 48560
rect 12820 48346 12848 48622
rect 12440 48340 12492 48346
rect 12440 48282 12492 48288
rect 12808 48340 12860 48346
rect 12808 48282 12860 48288
rect 14372 48068 14424 48074
rect 14372 48010 14424 48016
rect 14384 47802 14412 48010
rect 14372 47796 14424 47802
rect 14372 47738 14424 47744
rect 14280 47660 14332 47666
rect 14280 47602 14332 47608
rect 14292 47258 14320 47602
rect 13268 47252 13320 47258
rect 13268 47194 13320 47200
rect 14280 47252 14332 47258
rect 14280 47194 14332 47200
rect 12084 41386 12204 41414
rect 11612 35012 11664 35018
rect 11612 34954 11664 34960
rect 11624 34746 11652 34954
rect 11612 34740 11664 34746
rect 11612 34682 11664 34688
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 11980 34604 12032 34610
rect 11980 34546 12032 34552
rect 10968 32564 11020 32570
rect 10968 32506 11020 32512
rect 10876 32428 10928 32434
rect 10876 32370 10928 32376
rect 10888 32026 10916 32370
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 10980 31906 11008 32506
rect 10140 31884 10192 31890
rect 10140 31826 10192 31832
rect 10888 31878 11008 31906
rect 11244 31952 11296 31958
rect 11244 31894 11296 31900
rect 10152 30938 10180 31826
rect 10888 31822 10916 31878
rect 10876 31816 10928 31822
rect 10876 31758 10928 31764
rect 11152 31816 11204 31822
rect 11152 31758 11204 31764
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 8300 30660 8352 30666
rect 8300 30602 8352 30608
rect 8208 30320 8260 30326
rect 8208 30262 8260 30268
rect 8024 28484 8076 28490
rect 8024 28426 8076 28432
rect 8036 28218 8064 28426
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 8036 26994 8064 28154
rect 8220 28082 8248 30262
rect 8312 30258 8340 30602
rect 9956 30592 10008 30598
rect 9956 30534 10008 30540
rect 9680 30388 9732 30394
rect 9680 30330 9732 30336
rect 8300 30252 8352 30258
rect 8300 30194 8352 30200
rect 9312 30048 9364 30054
rect 9312 29990 9364 29996
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 8576 28484 8628 28490
rect 8576 28426 8628 28432
rect 8484 28416 8536 28422
rect 8484 28358 8536 28364
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8496 27470 8524 28358
rect 8588 27878 8616 28426
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8576 27872 8628 27878
rect 8576 27814 8628 27820
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8208 27328 8260 27334
rect 8208 27270 8260 27276
rect 8024 26988 8076 26994
rect 8024 26930 8076 26936
rect 8220 26926 8248 27270
rect 8208 26920 8260 26926
rect 8208 26862 8260 26868
rect 8588 26450 8616 27814
rect 8956 27606 8984 27950
rect 8944 27600 8996 27606
rect 8944 27542 8996 27548
rect 9140 27538 9168 28494
rect 9128 27532 9180 27538
rect 9128 27474 9180 27480
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 9128 26308 9180 26314
rect 9128 26250 9180 26256
rect 9140 26042 9168 26250
rect 9128 26036 9180 26042
rect 9128 25978 9180 25984
rect 8300 25900 8352 25906
rect 8300 25842 8352 25848
rect 8312 25226 8340 25842
rect 9232 25838 9260 29174
rect 9324 25906 9352 29990
rect 9692 29578 9720 30330
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9692 28914 9720 29514
rect 9968 29306 9996 30534
rect 10060 29646 10088 30670
rect 10048 29640 10100 29646
rect 10048 29582 10100 29588
rect 10060 29306 10088 29582
rect 10152 29510 10180 30874
rect 10416 30728 10468 30734
rect 10416 30670 10468 30676
rect 10428 30394 10456 30670
rect 10416 30388 10468 30394
rect 10416 30330 10468 30336
rect 10324 30252 10376 30258
rect 10324 30194 10376 30200
rect 10336 29850 10364 30194
rect 10324 29844 10376 29850
rect 10324 29786 10376 29792
rect 10600 29640 10652 29646
rect 10600 29582 10652 29588
rect 10140 29504 10192 29510
rect 10140 29446 10192 29452
rect 9956 29300 10008 29306
rect 9956 29242 10008 29248
rect 10048 29300 10100 29306
rect 10048 29242 10100 29248
rect 10060 29170 10088 29242
rect 10048 29164 10100 29170
rect 10048 29106 10100 29112
rect 9692 28886 9812 28914
rect 9496 28688 9548 28694
rect 9496 28630 9548 28636
rect 9404 28552 9456 28558
rect 9404 28494 9456 28500
rect 9416 27130 9444 28494
rect 9508 27402 9536 28630
rect 9588 28552 9640 28558
rect 9588 28494 9640 28500
rect 9600 27470 9628 28494
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9692 27538 9720 28018
rect 9680 27532 9732 27538
rect 9680 27474 9732 27480
rect 9588 27464 9640 27470
rect 9588 27406 9640 27412
rect 9496 27396 9548 27402
rect 9496 27338 9548 27344
rect 9600 27130 9628 27406
rect 9784 27334 9812 28886
rect 10048 28756 10100 28762
rect 10048 28698 10100 28704
rect 9772 27328 9824 27334
rect 9772 27270 9824 27276
rect 9404 27124 9456 27130
rect 9404 27066 9456 27072
rect 9588 27124 9640 27130
rect 9588 27066 9640 27072
rect 9312 25900 9364 25906
rect 9312 25842 9364 25848
rect 9220 25832 9272 25838
rect 9220 25774 9272 25780
rect 9232 25362 9260 25774
rect 9772 25424 9824 25430
rect 9416 25372 9772 25378
rect 9416 25366 9824 25372
rect 9220 25356 9272 25362
rect 9220 25298 9272 25304
rect 9416 25350 9812 25366
rect 9864 25356 9916 25362
rect 8760 25288 8812 25294
rect 8760 25230 8812 25236
rect 8300 25220 8352 25226
rect 8300 25162 8352 25168
rect 8392 24812 8444 24818
rect 8392 24754 8444 24760
rect 8404 24410 8432 24754
rect 8772 24750 8800 25230
rect 9128 25152 9180 25158
rect 9312 25152 9364 25158
rect 9180 25112 9312 25140
rect 9128 25094 9180 25100
rect 9312 25094 9364 25100
rect 9416 24886 9444 25350
rect 9864 25298 9916 25304
rect 9588 25288 9640 25294
rect 9588 25230 9640 25236
rect 9404 24880 9456 24886
rect 9404 24822 9456 24828
rect 9220 24812 9272 24818
rect 9220 24754 9272 24760
rect 9600 24800 9628 25230
rect 9677 24812 9729 24818
rect 9600 24772 9677 24800
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 9232 24614 9260 24754
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 7760 22066 7972 22094
rect 7012 22024 7064 22030
rect 7012 21966 7064 21972
rect 7472 21480 7524 21486
rect 7472 21422 7524 21428
rect 6460 20868 6512 20874
rect 6460 20810 6512 20816
rect 6472 20602 6500 20810
rect 6460 20596 6512 20602
rect 6460 20538 6512 20544
rect 7484 20534 7512 21422
rect 7472 20528 7524 20534
rect 7472 20470 7524 20476
rect 6368 20460 6420 20466
rect 6368 20402 6420 20408
rect 6380 20262 6408 20402
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6196 6886 6316 6914
rect 6196 4078 6224 6886
rect 6276 4616 6328 4622
rect 6276 4558 6328 4564
rect 6184 4072 6236 4078
rect 6184 4014 6236 4020
rect 5172 3936 5224 3942
rect 5172 3878 5224 3884
rect 5540 3936 5592 3942
rect 5540 3878 5592 3884
rect 5184 3602 5212 3878
rect 5552 3602 5580 3878
rect 5172 3596 5224 3602
rect 5172 3538 5224 3544
rect 5540 3596 5592 3602
rect 5540 3538 5592 3544
rect 5172 3460 5224 3466
rect 5172 3402 5224 3408
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 3976 2644 4028 2650
rect 3976 2586 4028 2592
rect 4068 2644 4120 2650
rect 4068 2586 4120 2592
rect 4080 2145 4108 2586
rect 4528 2440 4580 2446
rect 4528 2382 4580 2388
rect 4802 2408 4858 2417
rect 4066 2136 4122 2145
rect 4066 2071 4122 2080
rect 4540 800 4568 2382
rect 4802 2343 4858 2352
rect 4816 2310 4844 2343
rect 4804 2304 4856 2310
rect 4804 2246 4856 2252
rect 5184 800 5212 3402
rect 6288 3058 6316 4558
rect 6380 4146 6408 20198
rect 7760 18834 7788 22066
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7852 19786 7880 20470
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7748 18828 7800 18834
rect 7748 18770 7800 18776
rect 7104 18760 7156 18766
rect 7104 18702 7156 18708
rect 6828 18624 6880 18630
rect 6828 18566 6880 18572
rect 6840 18358 6868 18566
rect 6828 18352 6880 18358
rect 6828 18294 6880 18300
rect 7116 13326 7144 18702
rect 7852 18426 7880 19722
rect 7932 19304 7984 19310
rect 7932 19246 7984 19252
rect 7944 18970 7972 19246
rect 7932 18964 7984 18970
rect 7932 18906 7984 18912
rect 8036 18766 8064 23054
rect 8208 22024 8260 22030
rect 8208 21966 8260 21972
rect 8220 21690 8248 21966
rect 8208 21684 8260 21690
rect 8208 21626 8260 21632
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8220 20602 8248 20742
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8208 19712 8260 19718
rect 8208 19654 8260 19660
rect 8220 19310 8248 19654
rect 8208 19304 8260 19310
rect 8208 19246 8260 19252
rect 8300 18828 8352 18834
rect 8300 18770 8352 18776
rect 8024 18760 8076 18766
rect 8024 18702 8076 18708
rect 7840 18420 7892 18426
rect 7840 18362 7892 18368
rect 7852 18222 7880 18362
rect 7840 18216 7892 18222
rect 7840 18158 7892 18164
rect 7380 17604 7432 17610
rect 7380 17546 7432 17552
rect 7392 17270 7420 17546
rect 7380 17264 7432 17270
rect 7380 17206 7432 17212
rect 7852 17202 7880 18158
rect 8312 17882 8340 18770
rect 8680 18766 8708 24550
rect 9600 24274 9628 24772
rect 9677 24754 9729 24760
rect 9588 24268 9640 24274
rect 9588 24210 9640 24216
rect 9036 24200 9088 24206
rect 9036 24142 9088 24148
rect 9680 24200 9732 24206
rect 9680 24142 9732 24148
rect 9048 20942 9076 24142
rect 9496 23724 9548 23730
rect 9496 23666 9548 23672
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 9036 20936 9088 20942
rect 9036 20878 9088 20884
rect 8944 20800 8996 20806
rect 8944 20742 8996 20748
rect 8956 20466 8984 20742
rect 8944 20460 8996 20466
rect 8944 20402 8996 20408
rect 8668 18760 8720 18766
rect 8668 18702 8720 18708
rect 8944 18624 8996 18630
rect 8944 18566 8996 18572
rect 8956 18358 8984 18566
rect 8944 18352 8996 18358
rect 8944 18294 8996 18300
rect 8760 18080 8812 18086
rect 8760 18022 8812 18028
rect 8300 17876 8352 17882
rect 8300 17818 8352 17824
rect 7932 17672 7984 17678
rect 7932 17614 7984 17620
rect 7944 17338 7972 17614
rect 8772 17542 8800 18022
rect 8760 17536 8812 17542
rect 8760 17478 8812 17484
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 7932 17332 7984 17338
rect 7932 17274 7984 17280
rect 7840 17196 7892 17202
rect 7840 17138 7892 17144
rect 7104 13320 7156 13326
rect 7104 13262 7156 13268
rect 7196 4616 7248 4622
rect 7196 4558 7248 4564
rect 6368 4140 6420 4146
rect 6368 4082 6420 4088
rect 7012 4140 7064 4146
rect 7012 4082 7064 4088
rect 7024 3602 7052 4082
rect 7104 3936 7156 3942
rect 7104 3878 7156 3884
rect 7012 3596 7064 3602
rect 7012 3538 7064 3544
rect 6920 3460 6972 3466
rect 6920 3402 6972 3408
rect 6276 3052 6328 3058
rect 6276 2994 6328 3000
rect 6644 2984 6696 2990
rect 6472 2932 6644 2938
rect 6472 2926 6696 2932
rect 6472 2910 6684 2926
rect 5816 2848 5868 2854
rect 5816 2790 5868 2796
rect 5828 800 5856 2790
rect 6472 800 6500 2910
rect 6932 2514 6960 3402
rect 7116 2922 7144 3878
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 7024 2514 7052 2790
rect 7208 2582 7236 4558
rect 7944 4146 7972 17274
rect 8956 17202 8984 17478
rect 8944 17196 8996 17202
rect 8944 17138 8996 17144
rect 8024 16652 8076 16658
rect 8024 16594 8076 16600
rect 8036 4622 8064 16594
rect 8024 4616 8076 4622
rect 8024 4558 8076 4564
rect 7932 4140 7984 4146
rect 7932 4082 7984 4088
rect 7932 3936 7984 3942
rect 7932 3878 7984 3884
rect 7944 3670 7972 3878
rect 8036 3670 8064 4558
rect 8116 4480 8168 4486
rect 8116 4422 8168 4428
rect 8128 4214 8156 4422
rect 8116 4208 8168 4214
rect 8116 4150 8168 4156
rect 7932 3664 7984 3670
rect 7932 3606 7984 3612
rect 8024 3664 8076 3670
rect 8024 3606 8076 3612
rect 9036 3528 9088 3534
rect 9036 3470 9088 3476
rect 7748 2984 7800 2990
rect 7748 2926 7800 2932
rect 7196 2576 7248 2582
rect 7196 2518 7248 2524
rect 6920 2508 6972 2514
rect 6920 2450 6972 2456
rect 7012 2508 7064 2514
rect 7012 2450 7064 2456
rect 7472 2508 7524 2514
rect 7472 2450 7524 2456
rect 7116 870 7236 898
rect 7116 800 7144 870
rect 2778 776 2834 785
rect 2778 711 2834 720
rect 3238 0 3294 800
rect 3882 0 3938 800
rect 4526 0 4582 800
rect 5170 0 5226 800
rect 5814 0 5870 800
rect 6458 0 6514 800
rect 7102 0 7158 800
rect 7208 762 7236 870
rect 7484 762 7512 2450
rect 7760 800 7788 2926
rect 8392 2372 8444 2378
rect 8392 2314 8444 2320
rect 8404 800 8432 2314
rect 9048 800 9076 3470
rect 9140 2650 9168 23598
rect 9508 23322 9536 23666
rect 9588 23656 9640 23662
rect 9588 23598 9640 23604
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9220 21956 9272 21962
rect 9220 21898 9272 21904
rect 9232 20466 9260 21898
rect 9404 21616 9456 21622
rect 9324 21576 9404 21604
rect 9324 20939 9352 21576
rect 9404 21558 9456 21564
rect 9508 21554 9536 23258
rect 9600 23050 9628 23598
rect 9692 23322 9720 24142
rect 9876 23526 9904 25298
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9968 24410 9996 24754
rect 9956 24404 10008 24410
rect 9956 24346 10008 24352
rect 10060 24138 10088 28698
rect 10612 28558 10640 29582
rect 10888 29510 10916 31758
rect 11164 30734 11192 31758
rect 11256 30870 11284 31894
rect 11520 31816 11572 31822
rect 11520 31758 11572 31764
rect 11244 30864 11296 30870
rect 11244 30806 11296 30812
rect 11532 30734 11560 31758
rect 11796 30864 11848 30870
rect 11796 30806 11848 30812
rect 11152 30728 11204 30734
rect 11152 30670 11204 30676
rect 11520 30728 11572 30734
rect 11520 30670 11572 30676
rect 10968 30388 11020 30394
rect 10968 30330 11020 30336
rect 10980 29850 11008 30330
rect 11164 30258 11192 30670
rect 11152 30252 11204 30258
rect 11152 30194 11204 30200
rect 11428 30184 11480 30190
rect 11428 30126 11480 30132
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 11336 29640 11388 29646
rect 11336 29582 11388 29588
rect 10876 29504 10928 29510
rect 10876 29446 10928 29452
rect 10888 28762 10916 29446
rect 11244 28960 11296 28966
rect 11244 28902 11296 28908
rect 11150 28792 11206 28801
rect 10876 28756 10928 28762
rect 11150 28727 11206 28736
rect 10876 28698 10928 28704
rect 11164 28694 11192 28727
rect 11152 28688 11204 28694
rect 11152 28630 11204 28636
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 11152 28484 11204 28490
rect 11152 28426 11204 28432
rect 10600 28416 10652 28422
rect 10600 28358 10652 28364
rect 11060 28416 11112 28422
rect 11060 28358 11112 28364
rect 10612 28150 10640 28358
rect 10600 28144 10652 28150
rect 10600 28086 10652 28092
rect 10784 27396 10836 27402
rect 10784 27338 10836 27344
rect 10232 27328 10284 27334
rect 10232 27270 10284 27276
rect 10244 25906 10272 27270
rect 10796 26994 10824 27338
rect 11072 27334 11100 28358
rect 11164 27606 11192 28426
rect 11256 28014 11284 28902
rect 11348 28694 11376 29582
rect 11440 29578 11468 30126
rect 11808 29714 11836 30806
rect 11796 29708 11848 29714
rect 11796 29650 11848 29656
rect 11428 29572 11480 29578
rect 11428 29514 11480 29520
rect 11336 28688 11388 28694
rect 11336 28630 11388 28636
rect 11336 28552 11388 28558
rect 11440 28540 11468 29514
rect 11796 29300 11848 29306
rect 11796 29242 11848 29248
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11532 28540 11560 28630
rect 11388 28512 11560 28540
rect 11336 28494 11388 28500
rect 11244 28008 11296 28014
rect 11244 27950 11296 27956
rect 11152 27600 11204 27606
rect 11152 27542 11204 27548
rect 11244 27600 11296 27606
rect 11244 27542 11296 27548
rect 11256 27334 11284 27542
rect 11060 27328 11112 27334
rect 11060 27270 11112 27276
rect 11244 27328 11296 27334
rect 11244 27270 11296 27276
rect 10784 26988 10836 26994
rect 10784 26930 10836 26936
rect 10508 26444 10560 26450
rect 10508 26386 10560 26392
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10324 24744 10376 24750
rect 10324 24686 10376 24692
rect 10336 24274 10364 24686
rect 10416 24404 10468 24410
rect 10416 24346 10468 24352
rect 10324 24268 10376 24274
rect 10324 24210 10376 24216
rect 10048 24132 10100 24138
rect 10048 24074 10100 24080
rect 10428 23730 10456 24346
rect 10416 23724 10468 23730
rect 10416 23666 10468 23672
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9680 23316 9732 23322
rect 9680 23258 9732 23264
rect 9772 23316 9824 23322
rect 9772 23258 9824 23264
rect 9588 23044 9640 23050
rect 9588 22986 9640 22992
rect 9496 21548 9548 21554
rect 9496 21490 9548 21496
rect 9496 21412 9548 21418
rect 9496 21354 9548 21360
rect 9309 20933 9361 20939
rect 9309 20875 9361 20881
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9321 20816 9352 20875
rect 9220 20460 9272 20466
rect 9220 20402 9272 20408
rect 9232 17542 9260 20402
rect 9324 18970 9352 20816
rect 9416 20602 9444 20878
rect 9508 20806 9536 21354
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 9508 20482 9536 20742
rect 9416 20454 9536 20482
rect 9312 18964 9364 18970
rect 9312 18906 9364 18912
rect 9324 17814 9352 18906
rect 9416 18902 9444 20454
rect 9600 19904 9628 22986
rect 9784 22982 9812 23258
rect 10324 23248 10376 23254
rect 10324 23190 10376 23196
rect 10336 23118 10364 23190
rect 10428 23186 10456 23666
rect 10416 23180 10468 23186
rect 10416 23122 10468 23128
rect 10324 23112 10376 23118
rect 10322 23080 10324 23089
rect 10376 23080 10378 23089
rect 10322 23015 10378 23024
rect 9772 22976 9824 22982
rect 9772 22918 9824 22924
rect 10232 22024 10284 22030
rect 10232 21966 10284 21972
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9784 21554 9812 21830
rect 10244 21554 10272 21966
rect 9772 21548 9824 21554
rect 9772 21490 9824 21496
rect 10232 21548 10284 21554
rect 10232 21490 10284 21496
rect 9508 19876 9628 19904
rect 9404 18896 9456 18902
rect 9404 18838 9456 18844
rect 9312 17808 9364 17814
rect 9312 17750 9364 17756
rect 9508 17610 9536 19876
rect 10416 19712 10468 19718
rect 10416 19654 10468 19660
rect 10428 18766 10456 19654
rect 9588 18760 9640 18766
rect 9588 18702 9640 18708
rect 10416 18760 10468 18766
rect 10416 18702 10468 18708
rect 9600 18154 9628 18702
rect 9588 18148 9640 18154
rect 9588 18090 9640 18096
rect 9600 17678 9628 18090
rect 10428 17678 10456 18702
rect 9588 17672 9640 17678
rect 9588 17614 9640 17620
rect 10416 17672 10468 17678
rect 10416 17614 10468 17620
rect 9496 17604 9548 17610
rect 9496 17546 9548 17552
rect 9220 17536 9272 17542
rect 9220 17478 9272 17484
rect 9312 17332 9364 17338
rect 9312 17274 9364 17280
rect 9324 16998 9352 17274
rect 9312 16992 9364 16998
rect 9312 16934 9364 16940
rect 10232 4208 10284 4214
rect 10232 4150 10284 4156
rect 10244 3058 10272 4150
rect 10324 4004 10376 4010
rect 10324 3946 10376 3952
rect 9680 3052 9732 3058
rect 9680 2994 9732 3000
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 9128 2644 9180 2650
rect 9128 2586 9180 2592
rect 9692 800 9720 2994
rect 10336 800 10364 3946
rect 10520 3534 10548 26386
rect 10968 25696 11020 25702
rect 10968 25638 11020 25644
rect 10784 25424 10836 25430
rect 10784 25366 10836 25372
rect 10796 25294 10824 25366
rect 10784 25288 10836 25294
rect 10784 25230 10836 25236
rect 10876 25288 10928 25294
rect 10876 25230 10928 25236
rect 10888 24614 10916 25230
rect 10980 24886 11008 25638
rect 11348 25430 11376 28494
rect 11808 28014 11836 29242
rect 11888 28416 11940 28422
rect 11888 28358 11940 28364
rect 11704 28008 11756 28014
rect 11704 27950 11756 27956
rect 11796 28008 11848 28014
rect 11796 27950 11848 27956
rect 11612 25832 11664 25838
rect 11612 25774 11664 25780
rect 11336 25424 11388 25430
rect 11336 25366 11388 25372
rect 10968 24880 11020 24886
rect 10968 24822 11020 24828
rect 11624 24750 11652 25774
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 10876 24608 10928 24614
rect 10876 24550 10928 24556
rect 11716 23730 11744 27950
rect 11808 27402 11836 27950
rect 11900 27470 11928 28358
rect 11888 27464 11940 27470
rect 11888 27406 11940 27412
rect 11796 27396 11848 27402
rect 11796 27338 11848 27344
rect 11992 24954 12020 34546
rect 12072 28552 12124 28558
rect 12070 28520 12072 28529
rect 12124 28520 12126 28529
rect 12070 28455 12126 28464
rect 12072 25696 12124 25702
rect 12072 25638 12124 25644
rect 12084 25430 12112 25638
rect 12072 25424 12124 25430
rect 12072 25366 12124 25372
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11612 23656 11664 23662
rect 11612 23598 11664 23604
rect 11978 23624 12034 23633
rect 11624 23322 11652 23598
rect 11978 23559 11980 23568
rect 12032 23559 12034 23568
rect 11980 23530 12032 23536
rect 11612 23316 11664 23322
rect 11612 23258 11664 23264
rect 11612 21956 11664 21962
rect 11612 21898 11664 21904
rect 10600 21888 10652 21894
rect 10600 21830 10652 21836
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 10612 21010 10640 21830
rect 10600 21004 10652 21010
rect 10600 20946 10652 20952
rect 10784 20868 10836 20874
rect 10784 20810 10836 20816
rect 10796 20466 10824 20810
rect 10966 20496 11022 20505
rect 10600 20460 10652 20466
rect 10600 20402 10652 20408
rect 10784 20460 10836 20466
rect 10966 20431 10968 20440
rect 10784 20402 10836 20408
rect 11020 20431 11022 20440
rect 10968 20402 11020 20408
rect 10612 19786 10640 20402
rect 10796 20058 10824 20402
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 11164 19854 11192 20198
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 10600 19780 10652 19786
rect 10600 19722 10652 19728
rect 10612 18698 10640 19722
rect 10600 18692 10652 18698
rect 10600 18634 10652 18640
rect 10612 18358 10640 18634
rect 10600 18352 10652 18358
rect 10968 18352 11020 18358
rect 10600 18294 10652 18300
rect 10966 18320 10968 18329
rect 11020 18320 11022 18329
rect 10876 18284 10928 18290
rect 10966 18255 11022 18264
rect 10876 18226 10928 18232
rect 10888 17882 10916 18226
rect 10876 17876 10928 17882
rect 10876 17818 10928 17824
rect 10888 16658 10916 17818
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10784 15428 10836 15434
rect 10784 15370 10836 15376
rect 10796 15162 10824 15370
rect 10784 15156 10836 15162
rect 10784 15098 10836 15104
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10704 4078 10732 14962
rect 10692 4072 10744 4078
rect 10692 4014 10744 4020
rect 10508 3528 10560 3534
rect 10508 3470 10560 3476
rect 10968 2916 11020 2922
rect 10968 2858 11020 2864
rect 10600 2304 10652 2310
rect 10600 2246 10652 2252
rect 10612 1970 10640 2246
rect 10600 1964 10652 1970
rect 10600 1906 10652 1912
rect 10980 800 11008 2858
rect 7208 734 7512 762
rect 7746 0 7802 800
rect 8390 0 8446 800
rect 9034 0 9090 800
rect 9678 0 9734 800
rect 10322 0 10378 800
rect 10966 0 11022 800
rect 11256 762 11284 21830
rect 11624 21690 11652 21898
rect 11612 21684 11664 21690
rect 11612 21626 11664 21632
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11992 19961 12020 20402
rect 12072 20392 12124 20398
rect 12176 20380 12204 41386
rect 13280 35154 13308 47194
rect 13084 35148 13136 35154
rect 13084 35090 13136 35096
rect 13268 35148 13320 35154
rect 13268 35090 13320 35096
rect 13096 34202 13124 35090
rect 13084 34196 13136 34202
rect 13084 34138 13136 34144
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 13912 33040 13964 33046
rect 13912 32982 13964 32988
rect 13268 32972 13320 32978
rect 13268 32914 13320 32920
rect 13280 32570 13308 32914
rect 13820 32904 13872 32910
rect 13820 32846 13872 32852
rect 13268 32564 13320 32570
rect 13268 32506 13320 32512
rect 12716 32224 12768 32230
rect 12716 32166 12768 32172
rect 12728 31822 12756 32166
rect 13176 31952 13228 31958
rect 13176 31894 13228 31900
rect 12716 31816 12768 31822
rect 12716 31758 12768 31764
rect 12728 31210 12756 31758
rect 13084 31748 13136 31754
rect 13084 31690 13136 31696
rect 13096 31482 13124 31690
rect 13084 31476 13136 31482
rect 13084 31418 13136 31424
rect 12992 31408 13044 31414
rect 12990 31376 12992 31385
rect 13044 31376 13046 31385
rect 12990 31311 13046 31320
rect 12716 31204 12768 31210
rect 12716 31146 12768 31152
rect 12728 30326 12756 31146
rect 12716 30320 12768 30326
rect 12716 30262 12768 30268
rect 12728 29170 12756 30262
rect 13084 30048 13136 30054
rect 13084 29990 13136 29996
rect 13096 29238 13124 29990
rect 13084 29232 13136 29238
rect 13084 29174 13136 29180
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12624 29096 12676 29102
rect 12624 29038 12676 29044
rect 12636 28558 12664 29038
rect 12440 28552 12492 28558
rect 12440 28494 12492 28500
rect 12624 28552 12676 28558
rect 12624 28494 12676 28500
rect 12452 28218 12480 28494
rect 12440 28212 12492 28218
rect 12440 28154 12492 28160
rect 12636 26994 12664 28494
rect 13084 27600 13136 27606
rect 13084 27542 13136 27548
rect 13096 27130 13124 27542
rect 13084 27124 13136 27130
rect 13084 27066 13136 27072
rect 12624 26988 12676 26994
rect 12624 26930 12676 26936
rect 12714 25936 12770 25945
rect 12714 25871 12770 25880
rect 12728 25770 12756 25871
rect 12716 25764 12768 25770
rect 12716 25706 12768 25712
rect 12256 25696 12308 25702
rect 12256 25638 12308 25644
rect 12268 25294 12296 25638
rect 13188 25430 13216 31894
rect 13280 31482 13308 32506
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13360 31340 13412 31346
rect 13360 31282 13412 31288
rect 13372 30394 13400 31282
rect 13832 31278 13860 32846
rect 13924 32230 13952 32982
rect 14096 32768 14148 32774
rect 14096 32710 14148 32716
rect 14108 32502 14136 32710
rect 14096 32496 14148 32502
rect 14384 32450 14412 33458
rect 14464 32768 14516 32774
rect 14464 32710 14516 32716
rect 14096 32438 14148 32444
rect 14292 32434 14412 32450
rect 14280 32428 14412 32434
rect 14332 32422 14412 32428
rect 14280 32370 14332 32376
rect 14004 32360 14056 32366
rect 14004 32302 14056 32308
rect 13912 32224 13964 32230
rect 13912 32166 13964 32172
rect 13820 31272 13872 31278
rect 13820 31214 13872 31220
rect 13728 31136 13780 31142
rect 13728 31078 13780 31084
rect 13360 30388 13412 30394
rect 13360 30330 13412 30336
rect 13740 30122 13768 31078
rect 13832 30190 13860 31214
rect 13924 30734 13952 32166
rect 14016 31346 14044 32302
rect 14384 31890 14412 32422
rect 14372 31884 14424 31890
rect 14372 31826 14424 31832
rect 14096 31476 14148 31482
rect 14096 31418 14148 31424
rect 14108 31385 14136 31418
rect 14094 31376 14150 31385
rect 14004 31340 14056 31346
rect 14384 31346 14412 31826
rect 14094 31311 14150 31320
rect 14372 31340 14424 31346
rect 14004 31282 14056 31288
rect 14372 31282 14424 31288
rect 13912 30728 13964 30734
rect 13912 30670 13964 30676
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13728 30116 13780 30122
rect 13728 30058 13780 30064
rect 13740 29714 13768 30058
rect 13924 29714 13952 30670
rect 14016 30190 14044 31282
rect 14280 30728 14332 30734
rect 14384 30716 14412 31282
rect 14476 31142 14504 32710
rect 14660 31396 14688 49030
rect 14924 48544 14976 48550
rect 14924 48486 14976 48492
rect 14936 48210 14964 48486
rect 15028 48210 15056 51326
rect 15212 51326 15530 51354
rect 14924 48204 14976 48210
rect 14924 48146 14976 48152
rect 15016 48204 15068 48210
rect 15016 48146 15068 48152
rect 15212 34474 15240 51326
rect 15474 51200 15530 51326
rect 16118 51354 16174 52000
rect 16762 51354 16818 52000
rect 16118 51326 16528 51354
rect 16118 51200 16174 51326
rect 16500 49314 16528 51326
rect 16762 51326 17080 51354
rect 16762 51200 16818 51326
rect 16500 49298 16620 49314
rect 16500 49292 16632 49298
rect 16500 49286 16580 49292
rect 16580 49234 16632 49240
rect 17052 48686 17080 51326
rect 17406 51200 17462 52000
rect 18050 51200 18106 52000
rect 18694 51200 18750 52000
rect 19338 51354 19394 52000
rect 19982 51354 20038 52000
rect 19338 51326 19472 51354
rect 19338 51200 19394 51326
rect 17224 49156 17276 49162
rect 17224 49098 17276 49104
rect 16856 48680 16908 48686
rect 16856 48622 16908 48628
rect 17040 48680 17092 48686
rect 17040 48622 17092 48628
rect 16672 48000 16724 48006
rect 16672 47942 16724 47948
rect 16684 47666 16712 47942
rect 16868 47802 16896 48622
rect 17132 48000 17184 48006
rect 17132 47942 17184 47948
rect 16856 47796 16908 47802
rect 16856 47738 16908 47744
rect 16672 47660 16724 47666
rect 16672 47602 16724 47608
rect 16684 47569 16712 47602
rect 16670 47560 16726 47569
rect 16670 47495 16726 47504
rect 17144 47190 17172 47942
rect 17132 47184 17184 47190
rect 17132 47126 17184 47132
rect 17236 41414 17264 49098
rect 17420 48278 17448 51200
rect 17960 49224 18012 49230
rect 17960 49166 18012 49172
rect 17592 49088 17644 49094
rect 17592 49030 17644 49036
rect 17408 48272 17460 48278
rect 17408 48214 17460 48220
rect 17408 48068 17460 48074
rect 17408 48010 17460 48016
rect 17420 47802 17448 48010
rect 17408 47796 17460 47802
rect 17408 47738 17460 47744
rect 17406 47560 17462 47569
rect 17406 47495 17408 47504
rect 17460 47495 17462 47504
rect 17408 47466 17460 47472
rect 17144 41386 17264 41414
rect 17040 38276 17092 38282
rect 17040 38218 17092 38224
rect 16488 37256 16540 37262
rect 16488 37198 16540 37204
rect 15568 36168 15620 36174
rect 15568 36110 15620 36116
rect 15580 35630 15608 36110
rect 16500 35630 16528 37198
rect 17052 36174 17080 38218
rect 17144 37942 17172 41386
rect 17408 39364 17460 39370
rect 17408 39306 17460 39312
rect 17224 39296 17276 39302
rect 17224 39238 17276 39244
rect 17132 37936 17184 37942
rect 17132 37878 17184 37884
rect 17236 37194 17264 39238
rect 17420 39098 17448 39306
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 17604 38962 17632 49030
rect 17972 48210 18000 49166
rect 18064 48754 18092 51200
rect 19444 49230 19472 51326
rect 19982 51326 20116 51354
rect 19982 51200 20038 51326
rect 20088 49230 20116 51326
rect 20626 51200 20682 52000
rect 21270 51200 21326 52000
rect 21914 51354 21970 52000
rect 21652 51326 21970 51354
rect 19432 49224 19484 49230
rect 19432 49166 19484 49172
rect 20076 49224 20128 49230
rect 20076 49166 20128 49172
rect 20536 49156 20588 49162
rect 20536 49098 20588 49104
rect 20352 49088 20404 49094
rect 20352 49030 20404 49036
rect 19574 48988 19882 49008
rect 19574 48986 19580 48988
rect 19636 48986 19660 48988
rect 19716 48986 19740 48988
rect 19796 48986 19820 48988
rect 19876 48986 19882 48988
rect 19636 48934 19638 48986
rect 19818 48934 19820 48986
rect 19574 48932 19580 48934
rect 19636 48932 19660 48934
rect 19716 48932 19740 48934
rect 19796 48932 19820 48934
rect 19876 48932 19882 48934
rect 19574 48912 19882 48932
rect 18052 48748 18104 48754
rect 18052 48690 18104 48696
rect 18052 48544 18104 48550
rect 18052 48486 18104 48492
rect 17960 48204 18012 48210
rect 17960 48146 18012 48152
rect 17776 47660 17828 47666
rect 17776 47602 17828 47608
rect 17592 38956 17644 38962
rect 17592 38898 17644 38904
rect 17224 37188 17276 37194
rect 17224 37130 17276 37136
rect 17684 37188 17736 37194
rect 17684 37130 17736 37136
rect 17408 36848 17460 36854
rect 17408 36790 17460 36796
rect 17132 36644 17184 36650
rect 17132 36586 17184 36592
rect 17144 36378 17172 36586
rect 17132 36372 17184 36378
rect 17132 36314 17184 36320
rect 17040 36168 17092 36174
rect 16960 36128 17040 36156
rect 15568 35624 15620 35630
rect 15568 35566 15620 35572
rect 16488 35624 16540 35630
rect 16488 35566 16540 35572
rect 15580 35290 15608 35566
rect 15568 35284 15620 35290
rect 15568 35226 15620 35232
rect 15580 34610 15608 35226
rect 15568 34604 15620 34610
rect 15568 34546 15620 34552
rect 15200 34468 15252 34474
rect 15200 34410 15252 34416
rect 15580 33998 15608 34546
rect 16396 34468 16448 34474
rect 16396 34410 16448 34416
rect 16408 34134 16436 34410
rect 16396 34128 16448 34134
rect 16396 34070 16448 34076
rect 15568 33992 15620 33998
rect 15568 33934 15620 33940
rect 15476 33924 15528 33930
rect 15476 33866 15528 33872
rect 15488 33658 15516 33866
rect 15476 33652 15528 33658
rect 15476 33594 15528 33600
rect 15580 32978 15608 33934
rect 15568 32972 15620 32978
rect 15568 32914 15620 32920
rect 16960 32910 16988 36128
rect 17040 36110 17092 36116
rect 17420 35766 17448 36790
rect 17696 36378 17724 37130
rect 17684 36372 17736 36378
rect 17684 36314 17736 36320
rect 17684 36168 17736 36174
rect 17684 36110 17736 36116
rect 17408 35760 17460 35766
rect 17408 35702 17460 35708
rect 17132 35488 17184 35494
rect 17132 35430 17184 35436
rect 17144 33862 17172 35430
rect 17420 35086 17448 35702
rect 17696 35222 17724 36110
rect 17684 35216 17736 35222
rect 17684 35158 17736 35164
rect 17408 35080 17460 35086
rect 17408 35022 17460 35028
rect 17684 34944 17736 34950
rect 17684 34886 17736 34892
rect 17696 34678 17724 34886
rect 17684 34672 17736 34678
rect 17684 34614 17736 34620
rect 17500 33924 17552 33930
rect 17500 33866 17552 33872
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 17052 33590 17080 33798
rect 17040 33584 17092 33590
rect 17040 33526 17092 33532
rect 17512 33522 17540 33866
rect 17500 33516 17552 33522
rect 17500 33458 17552 33464
rect 17684 33516 17736 33522
rect 17684 33458 17736 33464
rect 17132 33448 17184 33454
rect 17132 33390 17184 33396
rect 14740 32904 14792 32910
rect 14740 32846 14792 32852
rect 16948 32904 17000 32910
rect 16948 32846 17000 32852
rect 14752 31686 14780 32846
rect 16672 32836 16724 32842
rect 16672 32778 16724 32784
rect 16684 32570 16712 32778
rect 16672 32564 16724 32570
rect 16672 32506 16724 32512
rect 16580 32428 16632 32434
rect 16580 32370 16632 32376
rect 14740 31680 14792 31686
rect 14740 31622 14792 31628
rect 14740 31408 14792 31414
rect 14660 31368 14740 31396
rect 14740 31350 14792 31356
rect 15108 31272 15160 31278
rect 15108 31214 15160 31220
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14332 30688 14412 30716
rect 14280 30670 14332 30676
rect 14004 30184 14056 30190
rect 14004 30126 14056 30132
rect 13728 29708 13780 29714
rect 13728 29650 13780 29656
rect 13912 29708 13964 29714
rect 13912 29650 13964 29656
rect 13924 28665 13952 29650
rect 13910 28656 13966 28665
rect 14016 28626 14044 30126
rect 14292 29578 14320 30670
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14384 30326 14412 30534
rect 14372 30320 14424 30326
rect 14372 30262 14424 30268
rect 14280 29572 14332 29578
rect 14280 29514 14332 29520
rect 14096 29028 14148 29034
rect 14096 28970 14148 28976
rect 13910 28591 13966 28600
rect 14004 28620 14056 28626
rect 13820 28144 13872 28150
rect 13820 28086 13872 28092
rect 13268 27328 13320 27334
rect 13268 27270 13320 27276
rect 13280 27130 13308 27270
rect 13268 27124 13320 27130
rect 13268 27066 13320 27072
rect 13280 26314 13308 27066
rect 13832 26994 13860 28086
rect 13820 26988 13872 26994
rect 13820 26930 13872 26936
rect 13832 26790 13860 26930
rect 13820 26784 13872 26790
rect 13820 26726 13872 26732
rect 13268 26308 13320 26314
rect 13268 26250 13320 26256
rect 13280 25906 13308 26250
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13176 25424 13228 25430
rect 13176 25366 13228 25372
rect 12992 25356 13044 25362
rect 12992 25298 13044 25304
rect 12256 25288 12308 25294
rect 12256 25230 12308 25236
rect 12900 24404 12952 24410
rect 12900 24346 12952 24352
rect 12532 24132 12584 24138
rect 12532 24074 12584 24080
rect 12544 23730 12572 24074
rect 12808 24064 12860 24070
rect 12808 24006 12860 24012
rect 12624 23860 12676 23866
rect 12624 23802 12676 23808
rect 12636 23746 12664 23802
rect 12532 23724 12584 23730
rect 12636 23718 12756 23746
rect 12820 23730 12848 24006
rect 12912 23866 12940 24346
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 12532 23666 12584 23672
rect 12624 23588 12676 23594
rect 12624 23530 12676 23536
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12544 23322 12572 23462
rect 12532 23316 12584 23322
rect 12532 23258 12584 23264
rect 12636 23186 12664 23530
rect 12728 23526 12756 23718
rect 12808 23724 12860 23730
rect 12808 23666 12860 23672
rect 12716 23520 12768 23526
rect 12716 23462 12768 23468
rect 12624 23180 12676 23186
rect 12624 23122 12676 23128
rect 12820 22710 12848 23666
rect 13004 23322 13032 25298
rect 13188 24818 13216 25366
rect 13176 24812 13228 24818
rect 13176 24754 13228 24760
rect 13280 24138 13308 25842
rect 13452 25356 13504 25362
rect 13452 25298 13504 25304
rect 13464 24614 13492 25298
rect 13924 25294 13952 28591
rect 14004 28562 14056 28568
rect 14108 26926 14136 28970
rect 14280 28620 14332 28626
rect 14280 28562 14332 28568
rect 14292 28218 14320 28562
rect 14384 28558 14412 30262
rect 14464 30252 14516 30258
rect 14464 30194 14516 30200
rect 14476 30054 14504 30194
rect 14464 30048 14516 30054
rect 14464 29990 14516 29996
rect 14476 29306 14504 29990
rect 14464 29300 14516 29306
rect 14464 29242 14516 29248
rect 14476 28626 14504 29242
rect 14740 28688 14792 28694
rect 14740 28630 14792 28636
rect 14464 28620 14516 28626
rect 14464 28562 14516 28568
rect 14752 28558 14780 28630
rect 14372 28552 14424 28558
rect 14372 28494 14424 28500
rect 14740 28552 14792 28558
rect 14740 28494 14792 28500
rect 14280 28212 14332 28218
rect 14280 28154 14332 28160
rect 14280 27328 14332 27334
rect 14280 27270 14332 27276
rect 14096 26920 14148 26926
rect 14096 26862 14148 26868
rect 14188 26920 14240 26926
rect 14188 26862 14240 26868
rect 13912 25288 13964 25294
rect 13912 25230 13964 25236
rect 13544 25152 13596 25158
rect 13544 25094 13596 25100
rect 13452 24608 13504 24614
rect 13452 24550 13504 24556
rect 13268 24132 13320 24138
rect 13268 24074 13320 24080
rect 13084 24064 13136 24070
rect 13084 24006 13136 24012
rect 12992 23316 13044 23322
rect 12992 23258 13044 23264
rect 13096 23118 13124 24006
rect 13360 23724 13412 23730
rect 13360 23666 13412 23672
rect 13084 23112 13136 23118
rect 13084 23054 13136 23060
rect 12808 22704 12860 22710
rect 12808 22646 12860 22652
rect 13372 22642 13400 23666
rect 13268 22636 13320 22642
rect 13268 22578 13320 22584
rect 13360 22636 13412 22642
rect 13360 22578 13412 22584
rect 13176 22568 13228 22574
rect 13176 22510 13228 22516
rect 12992 22024 13044 22030
rect 13188 22012 13216 22510
rect 13280 22094 13308 22578
rect 13372 22234 13400 22578
rect 13464 22574 13492 24550
rect 13556 23662 13584 25094
rect 13728 23860 13780 23866
rect 13728 23802 13780 23808
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13636 22976 13688 22982
rect 13636 22918 13688 22924
rect 13648 22710 13676 22918
rect 13636 22704 13688 22710
rect 13636 22646 13688 22652
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13636 22568 13688 22574
rect 13636 22510 13688 22516
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13280 22066 13400 22094
rect 13188 21984 13308 22012
rect 12992 21966 13044 21972
rect 13004 21554 13032 21966
rect 13084 21956 13136 21962
rect 13084 21898 13136 21904
rect 12992 21548 13044 21554
rect 12992 21490 13044 21496
rect 13096 21350 13124 21898
rect 13084 21344 13136 21350
rect 13084 21286 13136 21292
rect 13176 20936 13228 20942
rect 13176 20878 13228 20884
rect 12438 20496 12494 20505
rect 12348 20460 12400 20466
rect 12438 20431 12440 20440
rect 12348 20402 12400 20408
rect 12492 20431 12494 20440
rect 12624 20460 12676 20466
rect 12440 20402 12492 20408
rect 12624 20402 12676 20408
rect 12124 20352 12204 20380
rect 12072 20334 12124 20340
rect 12256 20324 12308 20330
rect 12256 20266 12308 20272
rect 12268 20233 12296 20266
rect 12254 20224 12310 20233
rect 12254 20159 12310 20168
rect 12256 19984 12308 19990
rect 11978 19952 12034 19961
rect 12256 19926 12308 19932
rect 11978 19887 12034 19896
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 11796 19848 11848 19854
rect 11796 19790 11848 19796
rect 11808 19514 11836 19790
rect 11978 19544 12034 19553
rect 11796 19508 11848 19514
rect 11978 19479 12034 19488
rect 11796 19450 11848 19456
rect 11808 18970 11836 19450
rect 11992 19378 12020 19479
rect 11980 19372 12032 19378
rect 11980 19314 12032 19320
rect 12084 19258 12112 19858
rect 12164 19440 12216 19446
rect 12268 19428 12296 19926
rect 12360 19922 12388 20402
rect 12348 19916 12400 19922
rect 12400 19876 12480 19904
rect 12348 19858 12400 19864
rect 12452 19514 12480 19876
rect 12636 19825 12664 20402
rect 12992 19848 13044 19854
rect 12622 19816 12678 19825
rect 12992 19790 13044 19796
rect 12622 19751 12678 19760
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12216 19400 12296 19428
rect 12164 19382 12216 19388
rect 11900 19230 12112 19258
rect 11796 18964 11848 18970
rect 11796 18906 11848 18912
rect 11900 18850 11928 19230
rect 12072 19168 12124 19174
rect 12072 19110 12124 19116
rect 11980 18964 12032 18970
rect 11980 18906 12032 18912
rect 11808 18822 11928 18850
rect 11808 18222 11836 18822
rect 11888 18624 11940 18630
rect 11888 18566 11940 18572
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11900 18086 11928 18566
rect 11992 18290 12020 18906
rect 12084 18766 12112 19110
rect 12268 18834 12296 19400
rect 12636 19360 12664 19751
rect 12808 19712 12860 19718
rect 12808 19654 12860 19660
rect 12820 19446 12848 19654
rect 12808 19440 12860 19446
rect 12808 19382 12860 19388
rect 12716 19372 12768 19378
rect 12636 19332 12716 19360
rect 12716 19314 12768 19320
rect 12900 19236 12952 19242
rect 12900 19178 12952 19184
rect 12256 18828 12308 18834
rect 12256 18770 12308 18776
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12440 18760 12492 18766
rect 12440 18702 12492 18708
rect 12254 18320 12310 18329
rect 11980 18284 12032 18290
rect 12452 18290 12480 18702
rect 12912 18290 12940 19178
rect 12254 18255 12256 18264
rect 11980 18226 12032 18232
rect 12308 18255 12310 18264
rect 12440 18284 12492 18290
rect 12256 18226 12308 18232
rect 12440 18226 12492 18232
rect 12900 18284 12952 18290
rect 12900 18226 12952 18232
rect 11796 18080 11848 18086
rect 11796 18022 11848 18028
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 12900 18080 12952 18086
rect 12900 18022 12952 18028
rect 11808 17678 11836 18022
rect 11796 17672 11848 17678
rect 11796 17614 11848 17620
rect 11428 16652 11480 16658
rect 11428 16594 11480 16600
rect 11440 16454 11468 16594
rect 11612 16516 11664 16522
rect 11612 16458 11664 16464
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11624 16250 11652 16458
rect 11612 16244 11664 16250
rect 11612 16186 11664 16192
rect 11520 16108 11572 16114
rect 11520 16050 11572 16056
rect 11532 11762 11560 16050
rect 12348 15564 12400 15570
rect 12348 15506 12400 15512
rect 11520 11756 11572 11762
rect 11520 11698 11572 11704
rect 12360 4010 12388 15506
rect 12912 15502 12940 18022
rect 13004 17678 13032 19790
rect 13188 19378 13216 20878
rect 13280 19553 13308 21984
rect 13372 21554 13400 22066
rect 13648 21894 13676 22510
rect 13452 21888 13504 21894
rect 13452 21830 13504 21836
rect 13636 21888 13688 21894
rect 13636 21830 13688 21836
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 13372 19786 13400 21490
rect 13464 21350 13492 21830
rect 13740 21690 13768 23802
rect 14108 23050 14136 26862
rect 14200 25906 14228 26862
rect 14292 26858 14320 27270
rect 14384 27130 14412 28494
rect 14372 27124 14424 27130
rect 14372 27066 14424 27072
rect 14280 26852 14332 26858
rect 14280 26794 14332 26800
rect 14752 26518 14780 28494
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14844 27130 14872 27950
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 15016 27124 15068 27130
rect 15016 27066 15068 27072
rect 15028 26994 15056 27066
rect 15016 26988 15068 26994
rect 15016 26930 15068 26936
rect 14740 26512 14792 26518
rect 14740 26454 14792 26460
rect 14188 25900 14240 25906
rect 14188 25842 14240 25848
rect 14200 25294 14228 25842
rect 14280 25832 14332 25838
rect 14278 25800 14280 25809
rect 14332 25800 14334 25809
rect 14278 25735 14334 25744
rect 14464 25424 14516 25430
rect 14464 25366 14516 25372
rect 14476 25294 14504 25366
rect 14188 25288 14240 25294
rect 14188 25230 14240 25236
rect 14464 25288 14516 25294
rect 14464 25230 14516 25236
rect 14372 25152 14424 25158
rect 14372 25094 14424 25100
rect 14384 24750 14412 25094
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 15120 24614 15148 31214
rect 15212 30870 15240 31214
rect 15200 30864 15252 30870
rect 15200 30806 15252 30812
rect 16592 30258 16620 32370
rect 17144 32298 17172 33390
rect 17224 33312 17276 33318
rect 17224 33254 17276 33260
rect 17236 32434 17264 33254
rect 17224 32428 17276 32434
rect 17224 32370 17276 32376
rect 17132 32292 17184 32298
rect 17132 32234 17184 32240
rect 16764 31340 16816 31346
rect 16764 31282 16816 31288
rect 16580 30252 16632 30258
rect 16580 30194 16632 30200
rect 16776 30122 16804 31282
rect 16856 30932 16908 30938
rect 16856 30874 16908 30880
rect 16580 30116 16632 30122
rect 16580 30058 16632 30064
rect 16764 30116 16816 30122
rect 16764 30058 16816 30064
rect 16592 30002 16620 30058
rect 16592 29974 16804 30002
rect 15844 29572 15896 29578
rect 15844 29514 15896 29520
rect 16028 29572 16080 29578
rect 16028 29514 16080 29520
rect 15292 29504 15344 29510
rect 15292 29446 15344 29452
rect 15304 29306 15332 29446
rect 15292 29300 15344 29306
rect 15292 29242 15344 29248
rect 15660 29096 15712 29102
rect 15660 29038 15712 29044
rect 15672 28801 15700 29038
rect 15658 28792 15714 28801
rect 15658 28727 15714 28736
rect 15856 28626 15884 29514
rect 15936 29504 15988 29510
rect 15936 29446 15988 29452
rect 15948 29170 15976 29446
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 16040 29073 16068 29514
rect 16304 29504 16356 29510
rect 16304 29446 16356 29452
rect 16316 29170 16344 29446
rect 16488 29232 16540 29238
rect 16488 29174 16540 29180
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 16026 29064 16082 29073
rect 16026 28999 16082 29008
rect 15844 28620 15896 28626
rect 15844 28562 15896 28568
rect 15856 28082 15884 28562
rect 15844 28076 15896 28082
rect 15844 28018 15896 28024
rect 16132 27606 16160 29106
rect 16500 28558 16528 29174
rect 16580 28960 16632 28966
rect 16580 28902 16632 28908
rect 16592 28626 16620 28902
rect 16776 28801 16804 29974
rect 16762 28792 16818 28801
rect 16762 28727 16818 28736
rect 16580 28620 16632 28626
rect 16580 28562 16632 28568
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16776 28218 16804 28727
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 16672 27600 16724 27606
rect 16672 27542 16724 27548
rect 15752 27532 15804 27538
rect 15752 27474 15804 27480
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 15660 27124 15712 27130
rect 15660 27066 15712 27072
rect 15672 26586 15700 27066
rect 15764 26994 15792 27474
rect 16396 27464 16448 27470
rect 16396 27406 16448 27412
rect 16304 27328 16356 27334
rect 16304 27270 16356 27276
rect 15752 26988 15804 26994
rect 15752 26930 15804 26936
rect 16316 26858 16344 27270
rect 16408 26926 16436 27406
rect 16396 26920 16448 26926
rect 16396 26862 16448 26868
rect 15752 26852 15804 26858
rect 15752 26794 15804 26800
rect 16304 26852 16356 26858
rect 16304 26794 16356 26800
rect 15764 26586 15792 26794
rect 15660 26580 15712 26586
rect 15660 26522 15712 26528
rect 15752 26580 15804 26586
rect 15752 26522 15804 26528
rect 16408 26382 16436 26862
rect 15384 26376 15436 26382
rect 16396 26376 16448 26382
rect 15384 26318 15436 26324
rect 15474 26344 15530 26353
rect 15396 25362 15424 26318
rect 16396 26318 16448 26324
rect 15474 26279 15476 26288
rect 15528 26279 15530 26288
rect 15476 26250 15528 26256
rect 16210 25664 16266 25673
rect 16210 25599 16266 25608
rect 16224 25362 16252 25599
rect 15384 25356 15436 25362
rect 15384 25298 15436 25304
rect 16212 25356 16264 25362
rect 16212 25298 16264 25304
rect 16592 25158 16620 27474
rect 16684 26994 16712 27542
rect 16672 26988 16724 26994
rect 16672 26930 16724 26936
rect 16684 26586 16712 26930
rect 16764 26784 16816 26790
rect 16764 26726 16816 26732
rect 16672 26580 16724 26586
rect 16672 26522 16724 26528
rect 16672 26308 16724 26314
rect 16672 26250 16724 26256
rect 16684 26042 16712 26250
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16776 25294 16804 26726
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 16580 25152 16632 25158
rect 16580 25094 16632 25100
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 14280 24608 14332 24614
rect 14280 24550 14332 24556
rect 15108 24608 15160 24614
rect 15108 24550 15160 24556
rect 14292 23798 14320 24550
rect 16592 24138 16620 24754
rect 16580 24132 16632 24138
rect 16580 24074 16632 24080
rect 14280 23792 14332 23798
rect 14280 23734 14332 23740
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14464 23520 14516 23526
rect 14464 23462 14516 23468
rect 14476 23322 14504 23462
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14096 23044 14148 23050
rect 14096 22986 14148 22992
rect 14108 22642 14136 22986
rect 14292 22710 14320 23258
rect 14462 23080 14518 23089
rect 14372 23044 14424 23050
rect 14462 23015 14518 23024
rect 14372 22986 14424 22992
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14384 22642 14412 22986
rect 14476 22982 14504 23015
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14096 22636 14148 22642
rect 14096 22578 14148 22584
rect 14372 22636 14424 22642
rect 14372 22578 14424 22584
rect 14280 22228 14332 22234
rect 14280 22170 14332 22176
rect 14188 22024 14240 22030
rect 14188 21966 14240 21972
rect 13728 21684 13780 21690
rect 13728 21626 13780 21632
rect 13452 21344 13504 21350
rect 13452 21286 13504 21292
rect 14004 21344 14056 21350
rect 14004 21286 14056 21292
rect 14016 20466 14044 21286
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 14004 20460 14056 20466
rect 14004 20402 14056 20408
rect 13452 20256 13504 20262
rect 13452 20198 13504 20204
rect 13360 19780 13412 19786
rect 13360 19722 13412 19728
rect 13266 19544 13322 19553
rect 13372 19514 13400 19722
rect 13266 19479 13322 19488
rect 13360 19508 13412 19514
rect 13176 19372 13228 19378
rect 13176 19314 13228 19320
rect 13188 17814 13216 19314
rect 13280 18154 13308 19479
rect 13360 19450 13412 19456
rect 13372 18970 13400 19450
rect 13464 19378 13492 20198
rect 13832 20058 13860 20402
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13452 19372 13504 19378
rect 13452 19314 13504 19320
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13924 18154 13952 20266
rect 14200 18290 14228 21966
rect 14292 21486 14320 22170
rect 14476 22166 14504 22646
rect 14568 22506 14596 23666
rect 14740 23520 14792 23526
rect 14740 23462 14792 23468
rect 14752 23186 14780 23462
rect 16592 23254 16620 24074
rect 16672 23520 16724 23526
rect 16672 23462 16724 23468
rect 16580 23248 16632 23254
rect 16580 23190 16632 23196
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 16684 23118 16712 23462
rect 15568 23112 15620 23118
rect 15568 23054 15620 23060
rect 16672 23112 16724 23118
rect 16672 23054 16724 23060
rect 15580 22574 15608 23054
rect 15568 22568 15620 22574
rect 15568 22510 15620 22516
rect 14556 22500 14608 22506
rect 14556 22442 14608 22448
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 16868 22094 16896 30874
rect 16948 30592 17000 30598
rect 16948 30534 17000 30540
rect 16960 30258 16988 30534
rect 17040 30320 17092 30326
rect 17040 30262 17092 30268
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17052 26994 17080 30262
rect 17144 28994 17172 32234
rect 17224 31816 17276 31822
rect 17224 31758 17276 31764
rect 17236 30666 17264 31758
rect 17512 31754 17540 33458
rect 17696 33046 17724 33458
rect 17684 33040 17736 33046
rect 17684 32982 17736 32988
rect 17592 32496 17644 32502
rect 17592 32438 17644 32444
rect 17328 31726 17540 31754
rect 17224 30660 17276 30666
rect 17224 30602 17276 30608
rect 17328 29170 17356 31726
rect 17408 30728 17460 30734
rect 17408 30670 17460 30676
rect 17420 30190 17448 30670
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17316 29164 17368 29170
rect 17316 29106 17368 29112
rect 17144 28966 17264 28994
rect 17328 28966 17356 29106
rect 17236 28490 17264 28966
rect 17316 28960 17368 28966
rect 17316 28902 17368 28908
rect 17420 28762 17448 29582
rect 17316 28756 17368 28762
rect 17316 28698 17368 28704
rect 17408 28756 17460 28762
rect 17408 28698 17460 28704
rect 17224 28484 17276 28490
rect 17224 28426 17276 28432
rect 17132 28076 17184 28082
rect 17132 28018 17184 28024
rect 17144 27470 17172 28018
rect 17236 28014 17264 28426
rect 17224 28008 17276 28014
rect 17224 27950 17276 27956
rect 17236 27674 17264 27950
rect 17328 27946 17356 28698
rect 17316 27940 17368 27946
rect 17316 27882 17368 27888
rect 17224 27668 17276 27674
rect 17224 27610 17276 27616
rect 17328 27470 17356 27882
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17512 27062 17540 30194
rect 17604 28626 17632 32438
rect 17684 30592 17736 30598
rect 17684 30534 17736 30540
rect 17696 29782 17724 30534
rect 17684 29776 17736 29782
rect 17684 29718 17736 29724
rect 17592 28620 17644 28626
rect 17592 28562 17644 28568
rect 17682 28520 17738 28529
rect 17682 28455 17738 28464
rect 17696 28422 17724 28455
rect 17684 28416 17736 28422
rect 17684 28358 17736 28364
rect 17788 28200 17816 47602
rect 17868 38820 17920 38826
rect 17868 38762 17920 38768
rect 17880 38486 17908 38762
rect 17868 38480 17920 38486
rect 17868 38422 17920 38428
rect 17880 33590 17908 38422
rect 18064 36786 18092 48486
rect 20260 48068 20312 48074
rect 20260 48010 20312 48016
rect 19574 47900 19882 47920
rect 19574 47898 19580 47900
rect 19636 47898 19660 47900
rect 19716 47898 19740 47900
rect 19796 47898 19820 47900
rect 19876 47898 19882 47900
rect 19636 47846 19638 47898
rect 19818 47846 19820 47898
rect 19574 47844 19580 47846
rect 19636 47844 19660 47846
rect 19716 47844 19740 47846
rect 19796 47844 19820 47846
rect 19876 47844 19882 47846
rect 19574 47824 19882 47844
rect 20272 47802 20300 48010
rect 20260 47796 20312 47802
rect 20260 47738 20312 47744
rect 20168 47660 20220 47666
rect 20168 47602 20220 47608
rect 19574 46812 19882 46832
rect 19574 46810 19580 46812
rect 19636 46810 19660 46812
rect 19716 46810 19740 46812
rect 19796 46810 19820 46812
rect 19876 46810 19882 46812
rect 19636 46758 19638 46810
rect 19818 46758 19820 46810
rect 19574 46756 19580 46758
rect 19636 46756 19660 46758
rect 19716 46756 19740 46758
rect 19796 46756 19820 46758
rect 19876 46756 19882 46758
rect 19574 46736 19882 46756
rect 19574 45724 19882 45744
rect 19574 45722 19580 45724
rect 19636 45722 19660 45724
rect 19716 45722 19740 45724
rect 19796 45722 19820 45724
rect 19876 45722 19882 45724
rect 19636 45670 19638 45722
rect 19818 45670 19820 45722
rect 19574 45668 19580 45670
rect 19636 45668 19660 45670
rect 19716 45668 19740 45670
rect 19796 45668 19820 45670
rect 19876 45668 19882 45670
rect 19574 45648 19882 45668
rect 19574 44636 19882 44656
rect 19574 44634 19580 44636
rect 19636 44634 19660 44636
rect 19716 44634 19740 44636
rect 19796 44634 19820 44636
rect 19876 44634 19882 44636
rect 19636 44582 19638 44634
rect 19818 44582 19820 44634
rect 19574 44580 19580 44582
rect 19636 44580 19660 44582
rect 19716 44580 19740 44582
rect 19796 44580 19820 44582
rect 19876 44580 19882 44582
rect 19574 44560 19882 44580
rect 19574 43548 19882 43568
rect 19574 43546 19580 43548
rect 19636 43546 19660 43548
rect 19716 43546 19740 43548
rect 19796 43546 19820 43548
rect 19876 43546 19882 43548
rect 19636 43494 19638 43546
rect 19818 43494 19820 43546
rect 19574 43492 19580 43494
rect 19636 43492 19660 43494
rect 19716 43492 19740 43494
rect 19796 43492 19820 43494
rect 19876 43492 19882 43494
rect 19574 43472 19882 43492
rect 19574 42460 19882 42480
rect 19574 42458 19580 42460
rect 19636 42458 19660 42460
rect 19716 42458 19740 42460
rect 19796 42458 19820 42460
rect 19876 42458 19882 42460
rect 19636 42406 19638 42458
rect 19818 42406 19820 42458
rect 19574 42404 19580 42406
rect 19636 42404 19660 42406
rect 19716 42404 19740 42406
rect 19796 42404 19820 42406
rect 19876 42404 19882 42406
rect 19574 42384 19882 42404
rect 19340 41608 19392 41614
rect 19340 41550 19392 41556
rect 18788 41064 18840 41070
rect 18788 41006 18840 41012
rect 18604 40520 18656 40526
rect 18604 40462 18656 40468
rect 18512 40044 18564 40050
rect 18512 39986 18564 39992
rect 18524 38962 18552 39986
rect 18512 38956 18564 38962
rect 18512 38898 18564 38904
rect 18420 38412 18472 38418
rect 18420 38354 18472 38360
rect 18432 38214 18460 38354
rect 18524 38282 18552 38898
rect 18616 38706 18644 40462
rect 18800 39914 18828 41006
rect 19156 40044 19208 40050
rect 19156 39986 19208 39992
rect 18788 39908 18840 39914
rect 18788 39850 18840 39856
rect 18800 39302 18828 39850
rect 19168 39642 19196 39986
rect 19352 39846 19380 41550
rect 19432 41472 19484 41478
rect 19432 41414 19484 41420
rect 19444 41274 19472 41414
rect 19574 41372 19882 41392
rect 19574 41370 19580 41372
rect 19636 41370 19660 41372
rect 19716 41370 19740 41372
rect 19796 41370 19820 41372
rect 19876 41370 19882 41372
rect 19636 41318 19638 41370
rect 19818 41318 19820 41370
rect 19574 41316 19580 41318
rect 19636 41316 19660 41318
rect 19716 41316 19740 41318
rect 19796 41316 19820 41318
rect 19876 41316 19882 41318
rect 19574 41296 19882 41316
rect 19432 41268 19484 41274
rect 19432 41210 19484 41216
rect 20076 41132 20128 41138
rect 20076 41074 20128 41080
rect 19984 40928 20036 40934
rect 19984 40870 20036 40876
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19340 39840 19392 39846
rect 19340 39782 19392 39788
rect 19156 39636 19208 39642
rect 19156 39578 19208 39584
rect 19352 39438 19380 39782
rect 19444 39506 19472 40326
rect 19574 40284 19882 40304
rect 19574 40282 19580 40284
rect 19636 40282 19660 40284
rect 19716 40282 19740 40284
rect 19796 40282 19820 40284
rect 19876 40282 19882 40284
rect 19636 40230 19638 40282
rect 19818 40230 19820 40282
rect 19574 40228 19580 40230
rect 19636 40228 19660 40230
rect 19716 40228 19740 40230
rect 19796 40228 19820 40230
rect 19876 40228 19882 40230
rect 19574 40208 19882 40228
rect 19892 40112 19944 40118
rect 19892 40054 19944 40060
rect 19432 39500 19484 39506
rect 19432 39442 19484 39448
rect 19904 39438 19932 40054
rect 19340 39432 19392 39438
rect 19340 39374 19392 39380
rect 19892 39432 19944 39438
rect 19892 39374 19944 39380
rect 18696 39296 18748 39302
rect 18696 39238 18748 39244
rect 18788 39296 18840 39302
rect 18788 39238 18840 39244
rect 18708 38894 18736 39238
rect 19574 39196 19882 39216
rect 19574 39194 19580 39196
rect 19636 39194 19660 39196
rect 19716 39194 19740 39196
rect 19796 39194 19820 39196
rect 19876 39194 19882 39196
rect 19636 39142 19638 39194
rect 19818 39142 19820 39194
rect 19574 39140 19580 39142
rect 19636 39140 19660 39142
rect 19716 39140 19740 39142
rect 19796 39140 19820 39142
rect 19876 39140 19882 39142
rect 19574 39120 19882 39140
rect 19708 39024 19760 39030
rect 19708 38966 19760 38972
rect 18696 38888 18748 38894
rect 18696 38830 18748 38836
rect 18788 38752 18840 38758
rect 18616 38678 18736 38706
rect 18788 38694 18840 38700
rect 18512 38276 18564 38282
rect 18512 38218 18564 38224
rect 18420 38208 18472 38214
rect 18420 38150 18472 38156
rect 18328 37868 18380 37874
rect 18328 37810 18380 37816
rect 18340 37466 18368 37810
rect 18432 37652 18460 38150
rect 18604 37664 18656 37670
rect 18432 37624 18552 37652
rect 18328 37460 18380 37466
rect 18328 37402 18380 37408
rect 18052 36780 18104 36786
rect 18052 36722 18104 36728
rect 18236 36780 18288 36786
rect 18236 36722 18288 36728
rect 18052 36644 18104 36650
rect 18052 36586 18104 36592
rect 17960 35692 18012 35698
rect 17960 35634 18012 35640
rect 17972 33658 18000 35634
rect 18064 35086 18092 36586
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 18156 35698 18184 36518
rect 18248 36378 18276 36722
rect 18328 36712 18380 36718
rect 18328 36654 18380 36660
rect 18236 36372 18288 36378
rect 18236 36314 18288 36320
rect 18340 36174 18368 36654
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18340 35766 18368 36110
rect 18524 36038 18552 37624
rect 18604 37606 18656 37612
rect 18616 36242 18644 37606
rect 18604 36236 18656 36242
rect 18604 36178 18656 36184
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18328 35760 18380 35766
rect 18328 35702 18380 35708
rect 18144 35692 18196 35698
rect 18144 35634 18196 35640
rect 18340 35086 18368 35702
rect 18049 35080 18101 35086
rect 18049 35022 18101 35028
rect 18144 35080 18196 35086
rect 18144 35022 18196 35028
rect 18328 35080 18380 35086
rect 18328 35022 18380 35028
rect 18156 34202 18184 35022
rect 18144 34196 18196 34202
rect 18144 34138 18196 34144
rect 17960 33652 18012 33658
rect 17960 33594 18012 33600
rect 17868 33584 17920 33590
rect 17868 33526 17920 33532
rect 17880 32570 17908 33526
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17868 32428 17920 32434
rect 17868 32370 17920 32376
rect 17880 31822 17908 32370
rect 17972 31890 18000 33594
rect 18144 32904 18196 32910
rect 18144 32846 18196 32852
rect 18156 32502 18184 32846
rect 18144 32496 18196 32502
rect 18144 32438 18196 32444
rect 18052 32428 18104 32434
rect 18052 32370 18104 32376
rect 17960 31884 18012 31890
rect 17960 31826 18012 31832
rect 17868 31816 17920 31822
rect 17868 31758 17920 31764
rect 17880 30938 17908 31758
rect 18064 31754 18092 32370
rect 18708 31754 18736 38678
rect 17960 31748 18092 31754
rect 18012 31726 18092 31748
rect 17960 31690 18012 31696
rect 18064 31142 18092 31726
rect 18616 31726 18736 31754
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17868 30932 17920 30938
rect 17868 30874 17920 30880
rect 18064 30802 18092 31078
rect 18052 30796 18104 30802
rect 18052 30738 18104 30744
rect 18512 30388 18564 30394
rect 18512 30330 18564 30336
rect 18420 30184 18472 30190
rect 18420 30126 18472 30132
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18144 30048 18196 30054
rect 18144 29990 18196 29996
rect 18064 29646 18092 29990
rect 18156 29850 18184 29990
rect 18432 29850 18460 30126
rect 18524 29850 18552 30330
rect 18144 29844 18196 29850
rect 18144 29786 18196 29792
rect 18420 29844 18472 29850
rect 18420 29786 18472 29792
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18052 29640 18104 29646
rect 18052 29582 18104 29588
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17696 28172 17816 28200
rect 17500 27056 17552 27062
rect 17500 26998 17552 27004
rect 17040 26988 17092 26994
rect 16960 26948 17040 26976
rect 16960 25906 16988 26948
rect 17040 26930 17092 26936
rect 17408 26988 17460 26994
rect 17408 26930 17460 26936
rect 17420 26586 17448 26930
rect 17040 26580 17092 26586
rect 17040 26522 17092 26528
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17052 26042 17080 26522
rect 17512 26518 17540 26998
rect 17696 26518 17724 28172
rect 17880 27062 17908 29106
rect 18050 29064 18106 29073
rect 18050 28999 18052 29008
rect 18104 28999 18106 29008
rect 18052 28970 18104 28976
rect 18236 28756 18288 28762
rect 18236 28698 18288 28704
rect 18052 28688 18104 28694
rect 18052 28630 18104 28636
rect 18142 28656 18198 28665
rect 18064 28150 18092 28630
rect 18142 28591 18198 28600
rect 18156 28558 18184 28591
rect 18144 28552 18196 28558
rect 18144 28494 18196 28500
rect 18052 28144 18104 28150
rect 18052 28086 18104 28092
rect 18248 28082 18276 28698
rect 18512 28552 18564 28558
rect 18512 28494 18564 28500
rect 18236 28076 18288 28082
rect 18236 28018 18288 28024
rect 17868 27056 17920 27062
rect 17868 26998 17920 27004
rect 17500 26512 17552 26518
rect 17500 26454 17552 26460
rect 17684 26512 17736 26518
rect 17684 26454 17736 26460
rect 17132 26376 17184 26382
rect 17696 26353 17724 26454
rect 17132 26318 17184 26324
rect 17682 26344 17738 26353
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 17144 25906 17172 26318
rect 17682 26279 17738 26288
rect 18248 26246 18276 28018
rect 18524 27130 18552 28494
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18512 26852 18564 26858
rect 18512 26794 18564 26800
rect 18524 26586 18552 26794
rect 18512 26580 18564 26586
rect 18512 26522 18564 26528
rect 18616 26382 18644 31726
rect 18800 31346 18828 38694
rect 19720 38282 19748 38966
rect 19800 38956 19852 38962
rect 19996 38944 20024 40870
rect 20088 40118 20116 41074
rect 20076 40112 20128 40118
rect 20076 40054 20128 40060
rect 20076 39432 20128 39438
rect 20076 39374 20128 39380
rect 19852 38916 20024 38944
rect 19800 38898 19852 38904
rect 19340 38276 19392 38282
rect 19340 38218 19392 38224
rect 19708 38276 19760 38282
rect 19708 38218 19760 38224
rect 19156 37392 19208 37398
rect 19156 37334 19208 37340
rect 19064 37324 19116 37330
rect 19064 37266 19116 37272
rect 18972 35216 19024 35222
rect 18972 35158 19024 35164
rect 18788 31340 18840 31346
rect 18788 31282 18840 31288
rect 18696 29504 18748 29510
rect 18696 29446 18748 29452
rect 18708 27470 18736 29446
rect 18788 28552 18840 28558
rect 18788 28494 18840 28500
rect 18800 28014 18828 28494
rect 18788 28008 18840 28014
rect 18788 27950 18840 27956
rect 18696 27464 18748 27470
rect 18696 27406 18748 27412
rect 18788 26988 18840 26994
rect 18788 26930 18840 26936
rect 18800 26874 18828 26930
rect 18800 26858 18920 26874
rect 18800 26852 18932 26858
rect 18800 26846 18880 26852
rect 18880 26794 18932 26800
rect 18604 26376 18656 26382
rect 18604 26318 18656 26324
rect 17316 26240 17368 26246
rect 17316 26182 17368 26188
rect 18236 26240 18288 26246
rect 18236 26182 18288 26188
rect 16948 25900 17000 25906
rect 16948 25842 17000 25848
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 16960 25702 16988 25842
rect 17144 25809 17172 25842
rect 17130 25800 17186 25809
rect 17130 25735 17186 25744
rect 16948 25696 17000 25702
rect 16948 25638 17000 25644
rect 17328 25430 17356 26182
rect 17408 25968 17460 25974
rect 17406 25936 17408 25945
rect 17460 25936 17462 25945
rect 17406 25871 17462 25880
rect 18236 25832 18288 25838
rect 18236 25774 18288 25780
rect 18248 25702 18276 25774
rect 17408 25696 17460 25702
rect 18236 25696 18288 25702
rect 17408 25638 17460 25644
rect 18234 25664 18236 25673
rect 18288 25664 18290 25673
rect 17316 25424 17368 25430
rect 17316 25366 17368 25372
rect 17040 25288 17092 25294
rect 17040 25230 17092 25236
rect 16684 22066 16896 22094
rect 14372 22024 14424 22030
rect 14372 21966 14424 21972
rect 14384 21894 14412 21966
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 15844 21888 15896 21894
rect 15844 21830 15896 21836
rect 14280 21480 14332 21486
rect 14280 21422 14332 21428
rect 14292 19961 14320 21422
rect 15660 21412 15712 21418
rect 15660 21354 15712 21360
rect 15672 21078 15700 21354
rect 15660 21072 15712 21078
rect 15660 21014 15712 21020
rect 14556 20868 14608 20874
rect 14556 20810 14608 20816
rect 14568 20602 14596 20810
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 15856 20466 15884 21830
rect 16488 20868 16540 20874
rect 16488 20810 16540 20816
rect 16500 20754 16528 20810
rect 16500 20726 16620 20754
rect 14924 20460 14976 20466
rect 14924 20402 14976 20408
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 15844 20460 15896 20466
rect 15844 20402 15896 20408
rect 14936 20058 14964 20402
rect 14924 20052 14976 20058
rect 14924 19994 14976 20000
rect 14278 19952 14334 19961
rect 14278 19887 14334 19896
rect 14292 19854 14320 19887
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 15120 19514 15148 20402
rect 15936 20392 15988 20398
rect 15934 20360 15936 20369
rect 15988 20360 15990 20369
rect 15934 20295 15990 20304
rect 15948 19786 15976 20295
rect 16120 19916 16172 19922
rect 16120 19858 16172 19864
rect 15936 19780 15988 19786
rect 15936 19722 15988 19728
rect 15108 19508 15160 19514
rect 15108 19450 15160 19456
rect 15120 18358 15148 19450
rect 16132 19446 16160 19858
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16592 19378 16620 20726
rect 15844 19372 15896 19378
rect 15844 19314 15896 19320
rect 16580 19372 16632 19378
rect 16580 19314 16632 19320
rect 15660 18896 15712 18902
rect 15660 18838 15712 18844
rect 15672 18358 15700 18838
rect 15752 18760 15804 18766
rect 15752 18702 15804 18708
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 14188 18284 14240 18290
rect 14188 18226 14240 18232
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 13268 18148 13320 18154
rect 13268 18090 13320 18096
rect 13912 18148 13964 18154
rect 13912 18090 13964 18096
rect 14004 18148 14056 18154
rect 14004 18090 14056 18096
rect 13176 17808 13228 17814
rect 13176 17750 13228 17756
rect 12992 17672 13044 17678
rect 12992 17614 13044 17620
rect 13188 17134 13216 17750
rect 13280 17678 13308 18090
rect 13452 18080 13504 18086
rect 13452 18022 13504 18028
rect 13268 17672 13320 17678
rect 13268 17614 13320 17620
rect 13464 17202 13492 18022
rect 13924 17814 13952 18090
rect 14016 17882 14044 18090
rect 14004 17876 14056 17882
rect 14004 17818 14056 17824
rect 13912 17808 13964 17814
rect 13912 17750 13964 17756
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13176 17128 13228 17134
rect 13176 17070 13228 17076
rect 13188 16726 13216 17070
rect 13176 16720 13228 16726
rect 13176 16662 13228 16668
rect 13728 16720 13780 16726
rect 13728 16662 13780 16668
rect 13740 16114 13768 16662
rect 13924 16658 13952 17750
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 13912 16652 13964 16658
rect 13912 16594 13964 16600
rect 13728 16108 13780 16114
rect 13728 16050 13780 16056
rect 14384 15638 14412 17546
rect 14568 17066 14596 18226
rect 15016 17128 15068 17134
rect 15016 17070 15068 17076
rect 14556 17060 14608 17066
rect 14556 17002 14608 17008
rect 14832 17060 14884 17066
rect 14832 17002 14884 17008
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14372 15632 14424 15638
rect 14372 15574 14424 15580
rect 12900 15496 12952 15502
rect 12900 15438 12952 15444
rect 12624 15360 12676 15366
rect 12624 15302 12676 15308
rect 12636 9674 12664 15302
rect 14568 10674 14596 16526
rect 14844 16522 14872 17002
rect 14832 16516 14884 16522
rect 14832 16458 14884 16464
rect 15028 16114 15056 17070
rect 15120 17066 15148 18294
rect 15384 18080 15436 18086
rect 15384 18022 15436 18028
rect 15108 17060 15160 17066
rect 15108 17002 15160 17008
rect 15120 16590 15148 17002
rect 15396 16658 15424 18022
rect 15476 17536 15528 17542
rect 15476 17478 15528 17484
rect 15488 17202 15516 17478
rect 15672 17354 15700 18294
rect 15764 17678 15792 18702
rect 15856 18290 15884 19314
rect 15844 18284 15896 18290
rect 15844 18226 15896 18232
rect 15752 17672 15804 17678
rect 15752 17614 15804 17620
rect 15580 17326 15700 17354
rect 15580 17270 15608 17326
rect 15568 17264 15620 17270
rect 15568 17206 15620 17212
rect 15476 17196 15528 17202
rect 15476 17138 15528 17144
rect 15660 17196 15712 17202
rect 15660 17138 15712 17144
rect 15672 17066 15700 17138
rect 15660 17060 15712 17066
rect 15660 17002 15712 17008
rect 15384 16652 15436 16658
rect 15384 16594 15436 16600
rect 15108 16584 15160 16590
rect 15108 16526 15160 16532
rect 15016 16108 15068 16114
rect 15016 16050 15068 16056
rect 15108 15904 15160 15910
rect 15108 15846 15160 15852
rect 15120 15638 15148 15846
rect 15108 15632 15160 15638
rect 15108 15574 15160 15580
rect 15764 14890 15792 17614
rect 15752 14884 15804 14890
rect 15752 14826 15804 14832
rect 15856 12782 15884 18226
rect 16580 17128 16632 17134
rect 16580 17070 16632 17076
rect 16592 16454 16620 17070
rect 16580 16448 16632 16454
rect 16580 16390 16632 16396
rect 15844 12776 15896 12782
rect 15844 12718 15896 12724
rect 14556 10668 14608 10674
rect 14556 10610 14608 10616
rect 12636 9646 12756 9674
rect 12532 4140 12584 4146
rect 12532 4082 12584 4088
rect 12440 4072 12492 4078
rect 12438 4040 12440 4049
rect 12492 4040 12494 4049
rect 12348 4004 12400 4010
rect 12438 3975 12494 3984
rect 12348 3946 12400 3952
rect 12544 3942 12572 4082
rect 11888 3936 11940 3942
rect 11888 3878 11940 3884
rect 12532 3936 12584 3942
rect 12532 3878 12584 3884
rect 11704 3528 11756 3534
rect 11704 3470 11756 3476
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11532 2854 11560 3334
rect 11624 3194 11652 3334
rect 11612 3188 11664 3194
rect 11612 3130 11664 3136
rect 11716 3058 11744 3470
rect 11900 3466 11928 3878
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12452 3466 12480 3674
rect 11888 3460 11940 3466
rect 11888 3402 11940 3408
rect 12440 3460 12492 3466
rect 12440 3402 12492 3408
rect 11704 3052 11756 3058
rect 11704 2994 11756 3000
rect 12728 2990 12756 9646
rect 16684 8362 16712 22066
rect 16764 20800 16816 20806
rect 16764 20742 16816 20748
rect 16856 20800 16908 20806
rect 16856 20742 16908 20748
rect 16776 20602 16804 20742
rect 16764 20596 16816 20602
rect 16764 20538 16816 20544
rect 16764 20460 16816 20466
rect 16868 20448 16896 20742
rect 16816 20420 16896 20448
rect 16764 20402 16816 20408
rect 16868 19854 16896 20420
rect 16856 19848 16908 19854
rect 16856 19790 16908 19796
rect 16856 19712 16908 19718
rect 16856 19654 16908 19660
rect 16868 19378 16896 19654
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16764 17536 16816 17542
rect 16764 17478 16816 17484
rect 16776 17202 16804 17478
rect 16764 17196 16816 17202
rect 16764 17138 16816 17144
rect 16948 17196 17000 17202
rect 16948 17138 17000 17144
rect 16960 16794 16988 17138
rect 16948 16788 17000 16794
rect 16948 16730 17000 16736
rect 17052 13938 17080 25230
rect 17132 24064 17184 24070
rect 17132 24006 17184 24012
rect 17224 24064 17276 24070
rect 17224 24006 17276 24012
rect 17144 23730 17172 24006
rect 17236 23798 17264 24006
rect 17224 23792 17276 23798
rect 17224 23734 17276 23740
rect 17132 23724 17184 23730
rect 17132 23666 17184 23672
rect 17236 23662 17264 23734
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17236 22710 17264 23598
rect 17224 22704 17276 22710
rect 17224 22646 17276 22652
rect 17316 21412 17368 21418
rect 17316 21354 17368 21360
rect 17328 20466 17356 21354
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17328 19514 17356 20402
rect 17316 19508 17368 19514
rect 17316 19450 17368 19456
rect 17420 17354 17448 25638
rect 18234 25599 18290 25608
rect 18248 25573 18276 25599
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18892 24614 18920 24754
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17972 23798 18000 24074
rect 18512 23860 18564 23866
rect 18512 23802 18564 23808
rect 17960 23792 18012 23798
rect 17960 23734 18012 23740
rect 18050 23760 18106 23769
rect 17500 23724 17552 23730
rect 17500 23666 17552 23672
rect 17512 21350 17540 23666
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17696 22545 17724 23462
rect 17880 22710 17908 23462
rect 17972 23050 18000 23734
rect 18524 23730 18552 23802
rect 18050 23695 18052 23704
rect 18104 23695 18106 23704
rect 18328 23724 18380 23730
rect 18052 23666 18104 23672
rect 18328 23666 18380 23672
rect 18512 23724 18564 23730
rect 18512 23666 18564 23672
rect 18340 23254 18368 23666
rect 18420 23656 18472 23662
rect 18418 23624 18420 23633
rect 18472 23624 18474 23633
rect 18418 23559 18474 23568
rect 18328 23248 18380 23254
rect 18328 23190 18380 23196
rect 18788 23112 18840 23118
rect 18788 23054 18840 23060
rect 17960 23044 18012 23050
rect 17960 22986 18012 22992
rect 18052 23044 18104 23050
rect 18052 22986 18104 22992
rect 17868 22704 17920 22710
rect 17868 22646 17920 22652
rect 17682 22536 17738 22545
rect 17682 22471 17738 22480
rect 18064 22098 18092 22986
rect 18800 22506 18828 23054
rect 18788 22500 18840 22506
rect 18788 22442 18840 22448
rect 18696 22432 18748 22438
rect 18696 22374 18748 22380
rect 18052 22092 18104 22098
rect 18708 22094 18736 22374
rect 18708 22066 18920 22094
rect 18052 22034 18104 22040
rect 18892 22030 18920 22066
rect 18420 22024 18472 22030
rect 18420 21966 18472 21972
rect 18512 22024 18564 22030
rect 18512 21966 18564 21972
rect 18788 22024 18840 22030
rect 18788 21966 18840 21972
rect 18880 22024 18932 22030
rect 18880 21966 18932 21972
rect 17868 21548 17920 21554
rect 17868 21490 17920 21496
rect 17500 21344 17552 21350
rect 17500 21286 17552 21292
rect 17880 21010 17908 21490
rect 18432 21418 18460 21966
rect 18524 21690 18552 21966
rect 18512 21684 18564 21690
rect 18512 21626 18564 21632
rect 18420 21412 18472 21418
rect 18420 21354 18472 21360
rect 18696 21140 18748 21146
rect 18696 21082 18748 21088
rect 17868 21004 17920 21010
rect 17868 20946 17920 20952
rect 17684 20528 17736 20534
rect 17684 20470 17736 20476
rect 17500 20324 17552 20330
rect 17500 20266 17552 20272
rect 17512 20233 17540 20266
rect 17696 20262 17724 20470
rect 18052 20460 18104 20466
rect 18052 20402 18104 20408
rect 17684 20256 17736 20262
rect 17498 20224 17554 20233
rect 17684 20198 17736 20204
rect 17498 20159 17554 20168
rect 17696 20058 17724 20198
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 19848 17736 19854
rect 17682 19816 17684 19825
rect 17736 19816 17738 19825
rect 17500 19780 17552 19786
rect 17682 19751 17738 19760
rect 17500 19722 17552 19728
rect 17512 18970 17540 19722
rect 17592 19372 17644 19378
rect 17592 19314 17644 19320
rect 17500 18964 17552 18970
rect 17500 18906 17552 18912
rect 17604 18358 17632 19314
rect 18064 18834 18092 20402
rect 18328 20392 18380 20398
rect 18328 20334 18380 20340
rect 18602 20360 18658 20369
rect 18236 19848 18288 19854
rect 18236 19790 18288 19796
rect 18248 19553 18276 19790
rect 18234 19544 18290 19553
rect 18144 19508 18196 19514
rect 18234 19479 18290 19488
rect 18144 19450 18196 19456
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18156 18766 18184 19450
rect 18340 19258 18368 20334
rect 18602 20295 18658 20304
rect 18616 20262 18644 20295
rect 18512 20256 18564 20262
rect 18512 20198 18564 20204
rect 18604 20256 18656 20262
rect 18604 20198 18656 20204
rect 18524 19854 18552 20198
rect 18708 19854 18736 21082
rect 18800 20806 18828 21966
rect 18788 20800 18840 20806
rect 18788 20742 18840 20748
rect 18512 19848 18564 19854
rect 18696 19848 18748 19854
rect 18512 19790 18564 19796
rect 18694 19816 18696 19825
rect 18748 19816 18750 19825
rect 18694 19751 18750 19760
rect 18340 19230 18460 19258
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 17592 18352 17644 18358
rect 17592 18294 17644 18300
rect 17604 17814 17632 18294
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 17592 17808 17644 17814
rect 17592 17750 17644 17756
rect 17684 17604 17736 17610
rect 17684 17546 17736 17552
rect 17328 17326 17448 17354
rect 17328 16114 17356 17326
rect 17408 17196 17460 17202
rect 17408 17138 17460 17144
rect 17592 17196 17644 17202
rect 17592 17138 17644 17144
rect 17420 16114 17448 17138
rect 17604 16794 17632 17138
rect 17500 16788 17552 16794
rect 17500 16730 17552 16736
rect 17592 16788 17644 16794
rect 17592 16730 17644 16736
rect 17512 16250 17540 16730
rect 17604 16590 17632 16730
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17696 16522 17724 17546
rect 17684 16516 17736 16522
rect 17684 16458 17736 16464
rect 17500 16244 17552 16250
rect 17500 16186 17552 16192
rect 17316 16108 17368 16114
rect 17316 16050 17368 16056
rect 17408 16108 17460 16114
rect 17408 16050 17460 16056
rect 17132 15904 17184 15910
rect 17132 15846 17184 15852
rect 17144 15434 17172 15846
rect 17420 15706 17448 16050
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17408 15700 17460 15706
rect 17408 15642 17460 15648
rect 17880 15638 17908 15982
rect 17868 15632 17920 15638
rect 17868 15574 17920 15580
rect 17132 15428 17184 15434
rect 17132 15370 17184 15376
rect 17040 13932 17092 13938
rect 17040 13874 17092 13880
rect 17316 13864 17368 13870
rect 17316 13806 17368 13812
rect 17328 13530 17356 13806
rect 17316 13524 17368 13530
rect 17316 13466 17368 13472
rect 16856 13320 16908 13326
rect 16856 13262 16908 13268
rect 16868 12850 16896 13262
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16948 12640 17000 12646
rect 16948 12582 17000 12588
rect 16960 11830 16988 12582
rect 16948 11824 17000 11830
rect 16948 11766 17000 11772
rect 16764 11688 16816 11694
rect 16764 11630 16816 11636
rect 16776 11354 16804 11630
rect 16764 11348 16816 11354
rect 16764 11290 16816 11296
rect 17316 11144 17368 11150
rect 17316 11086 17368 11092
rect 17328 9586 17356 11086
rect 17316 9580 17368 9586
rect 17316 9522 17368 9528
rect 17328 9042 17356 9522
rect 17316 9036 17368 9042
rect 17316 8978 17368 8984
rect 16672 8356 16724 8362
rect 16672 8298 16724 8304
rect 16488 7948 16540 7954
rect 16488 7890 16540 7896
rect 15200 6724 15252 6730
rect 15200 6666 15252 6672
rect 14924 4140 14976 4146
rect 14924 4082 14976 4088
rect 13176 4072 13228 4078
rect 13176 4014 13228 4020
rect 13544 4072 13596 4078
rect 13544 4014 13596 4020
rect 12808 3596 12860 3602
rect 12808 3538 12860 3544
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 12716 2984 12768 2990
rect 12716 2926 12768 2932
rect 11520 2848 11572 2854
rect 11520 2790 11572 2796
rect 12452 2650 12480 2926
rect 12440 2644 12492 2650
rect 12440 2586 12492 2592
rect 12820 1290 12848 3538
rect 12900 2984 12952 2990
rect 12900 2926 12952 2932
rect 12256 1284 12308 1290
rect 12256 1226 12308 1232
rect 12808 1284 12860 1290
rect 12808 1226 12860 1232
rect 11532 870 11652 898
rect 11532 762 11560 870
rect 11624 800 11652 870
rect 12268 800 12296 1226
rect 12912 800 12940 2926
rect 13188 2650 13216 4014
rect 13176 2644 13228 2650
rect 13176 2586 13228 2592
rect 13556 800 13584 4014
rect 14936 3534 14964 4082
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15120 3058 15148 3470
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 15212 2514 15240 6666
rect 15476 3392 15528 3398
rect 15476 3334 15528 3340
rect 15200 2508 15252 2514
rect 15200 2450 15252 2456
rect 14188 2372 14240 2378
rect 14188 2314 14240 2320
rect 14200 800 14228 2314
rect 15488 800 15516 3334
rect 16500 3126 16528 7890
rect 17972 4214 18000 18226
rect 18432 18154 18460 19230
rect 18800 18290 18828 20742
rect 18788 18284 18840 18290
rect 18788 18226 18840 18232
rect 18420 18148 18472 18154
rect 18420 18090 18472 18096
rect 18144 18080 18196 18086
rect 18144 18022 18196 18028
rect 18156 17202 18184 18022
rect 18236 17672 18288 17678
rect 18288 17632 18368 17660
rect 18236 17614 18288 17620
rect 18144 17196 18196 17202
rect 18144 17138 18196 17144
rect 18236 14884 18288 14890
rect 18236 14826 18288 14832
rect 18052 13864 18104 13870
rect 18052 13806 18104 13812
rect 18064 9722 18092 13806
rect 18248 12850 18276 14826
rect 18236 12844 18288 12850
rect 18236 12786 18288 12792
rect 18144 11688 18196 11694
rect 18144 11630 18196 11636
rect 18052 9716 18104 9722
rect 18052 9658 18104 9664
rect 17960 4208 18012 4214
rect 17960 4150 18012 4156
rect 17224 4072 17276 4078
rect 17224 4014 17276 4020
rect 17682 4040 17738 4049
rect 17236 3738 17264 4014
rect 17682 3975 17738 3984
rect 17316 3936 17368 3942
rect 17316 3878 17368 3884
rect 17224 3732 17276 3738
rect 17224 3674 17276 3680
rect 16488 3120 16540 3126
rect 16488 3062 16540 3068
rect 17328 3058 17356 3878
rect 17592 3732 17644 3738
rect 17592 3674 17644 3680
rect 17500 3392 17552 3398
rect 17500 3334 17552 3340
rect 17512 3126 17540 3334
rect 17500 3120 17552 3126
rect 17500 3062 17552 3068
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 17604 2990 17632 3674
rect 17696 3126 17724 3975
rect 17684 3120 17736 3126
rect 17684 3062 17736 3068
rect 17592 2984 17644 2990
rect 17592 2926 17644 2932
rect 18052 2984 18104 2990
rect 18052 2926 18104 2932
rect 17408 2372 17460 2378
rect 17408 2314 17460 2320
rect 17420 800 17448 2314
rect 18064 800 18092 2926
rect 18156 2854 18184 11630
rect 18340 3602 18368 17632
rect 18432 17542 18460 18090
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18512 17808 18564 17814
rect 18512 17750 18564 17756
rect 18524 17542 18552 17750
rect 18616 17610 18644 18022
rect 18800 17610 18828 18226
rect 18604 17604 18656 17610
rect 18604 17546 18656 17552
rect 18788 17604 18840 17610
rect 18788 17546 18840 17552
rect 18420 17536 18472 17542
rect 18420 17478 18472 17484
rect 18512 17536 18564 17542
rect 18512 17478 18564 17484
rect 18604 17332 18656 17338
rect 18604 17274 18656 17280
rect 18420 17264 18472 17270
rect 18616 17218 18644 17274
rect 18472 17212 18644 17218
rect 18420 17206 18644 17212
rect 18432 17190 18644 17206
rect 18420 16992 18472 16998
rect 18420 16934 18472 16940
rect 18788 16992 18840 16998
rect 18788 16934 18840 16940
rect 18432 16250 18460 16934
rect 18800 16726 18828 16934
rect 18788 16720 18840 16726
rect 18788 16662 18840 16668
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18708 14414 18736 16458
rect 18788 16108 18840 16114
rect 18788 16050 18840 16056
rect 18800 15434 18828 16050
rect 18788 15428 18840 15434
rect 18788 15370 18840 15376
rect 18696 14408 18748 14414
rect 18696 14350 18748 14356
rect 18880 8832 18932 8838
rect 18880 8774 18932 8780
rect 18696 8424 18748 8430
rect 18696 8366 18748 8372
rect 18708 8090 18736 8366
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18892 7886 18920 8774
rect 18880 7880 18932 7886
rect 18880 7822 18932 7828
rect 18892 7410 18920 7822
rect 18984 7750 19012 35158
rect 19076 32756 19104 37266
rect 19168 32910 19196 37334
rect 19352 37330 19380 38218
rect 19812 38196 19840 38898
rect 20088 38486 20116 39374
rect 20076 38480 20128 38486
rect 20076 38422 20128 38428
rect 19812 38168 20116 38196
rect 19574 38108 19882 38128
rect 19574 38106 19580 38108
rect 19636 38106 19660 38108
rect 19716 38106 19740 38108
rect 19796 38106 19820 38108
rect 19876 38106 19882 38108
rect 19636 38054 19638 38106
rect 19818 38054 19820 38106
rect 19574 38052 19580 38054
rect 19636 38052 19660 38054
rect 19716 38052 19740 38054
rect 19796 38052 19820 38054
rect 19876 38052 19882 38054
rect 19574 38032 19882 38052
rect 19432 37868 19484 37874
rect 19432 37810 19484 37816
rect 19340 37324 19392 37330
rect 19340 37266 19392 37272
rect 19340 36780 19392 36786
rect 19340 36722 19392 36728
rect 19248 36576 19300 36582
rect 19248 36518 19300 36524
rect 19260 36174 19288 36518
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19352 35494 19380 36722
rect 19444 36174 19472 37810
rect 19984 37324 20036 37330
rect 19984 37266 20036 37272
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19996 36904 20024 37266
rect 19904 36876 20024 36904
rect 19904 36718 19932 36876
rect 19892 36712 19944 36718
rect 19892 36654 19944 36660
rect 19904 36378 19932 36654
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19432 36168 19484 36174
rect 19432 36110 19484 36116
rect 19904 36122 19932 36314
rect 20088 36310 20116 38168
rect 20076 36304 20128 36310
rect 20076 36246 20128 36252
rect 19340 35488 19392 35494
rect 19340 35430 19392 35436
rect 19340 35080 19392 35086
rect 19340 35022 19392 35028
rect 19248 34944 19300 34950
rect 19248 34886 19300 34892
rect 19260 33998 19288 34886
rect 19352 34746 19380 35022
rect 19444 34746 19472 36110
rect 19904 36094 20024 36122
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19892 35760 19944 35766
rect 19892 35702 19944 35708
rect 19800 35488 19852 35494
rect 19798 35456 19800 35465
rect 19852 35456 19854 35465
rect 19798 35391 19854 35400
rect 19614 35184 19670 35193
rect 19614 35119 19670 35128
rect 19628 35086 19656 35119
rect 19616 35080 19668 35086
rect 19904 35057 19932 35702
rect 19996 35154 20024 36094
rect 20076 36032 20128 36038
rect 20076 35974 20128 35980
rect 19984 35148 20036 35154
rect 19984 35090 20036 35096
rect 19616 35022 19668 35028
rect 19890 35048 19946 35057
rect 19890 34983 19946 34992
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 19432 34740 19484 34746
rect 19432 34682 19484 34688
rect 19340 34604 19392 34610
rect 19340 34546 19392 34552
rect 19248 33992 19300 33998
rect 19248 33934 19300 33940
rect 19352 33522 19380 34546
rect 19444 33930 19472 34682
rect 19432 33924 19484 33930
rect 19432 33866 19484 33872
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19340 33516 19392 33522
rect 19340 33458 19392 33464
rect 19156 32904 19208 32910
rect 19156 32846 19208 32852
rect 19076 32728 19288 32756
rect 19260 31770 19288 32728
rect 19352 31890 19380 33458
rect 19432 32836 19484 32842
rect 19432 32778 19484 32784
rect 19340 31884 19392 31890
rect 19340 31826 19392 31832
rect 19260 31742 19380 31770
rect 19444 31754 19472 32778
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 19996 32450 20024 32710
rect 19904 32434 20024 32450
rect 19892 32428 20024 32434
rect 19944 32422 20024 32428
rect 19892 32370 19944 32376
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19260 31142 19288 31282
rect 19248 31136 19300 31142
rect 19248 31078 19300 31084
rect 19260 29714 19288 31078
rect 19248 29708 19300 29714
rect 19248 29650 19300 29656
rect 19352 29578 19380 31742
rect 19432 31748 19484 31754
rect 19432 31690 19484 31696
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19444 30258 19472 30534
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19432 30252 19484 30258
rect 19432 30194 19484 30200
rect 19444 29646 19472 30194
rect 19432 29640 19484 29646
rect 19432 29582 19484 29588
rect 19340 29572 19392 29578
rect 19340 29514 19392 29520
rect 19444 29238 19472 29582
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19522 29200 19578 29209
rect 19340 28960 19392 28966
rect 19340 28902 19392 28908
rect 19352 28098 19380 28902
rect 19444 28626 19472 29174
rect 19522 29135 19578 29144
rect 19432 28620 19484 28626
rect 19432 28562 19484 28568
rect 19168 28082 19380 28098
rect 19156 28076 19380 28082
rect 19208 28070 19380 28076
rect 19156 28018 19208 28024
rect 19444 27878 19472 28562
rect 19536 28404 19564 29135
rect 20088 28762 20116 35974
rect 20180 33017 20208 47602
rect 20364 47138 20392 49030
rect 20444 48544 20496 48550
rect 20444 48486 20496 48492
rect 20456 48210 20484 48486
rect 20444 48204 20496 48210
rect 20444 48146 20496 48152
rect 20548 47546 20576 49098
rect 20640 48210 20668 51200
rect 21652 49230 21680 51326
rect 21914 51200 21970 51326
rect 22558 51200 22614 52000
rect 23202 51354 23258 52000
rect 23202 51326 23428 51354
rect 23202 51200 23258 51326
rect 22572 49298 22600 51200
rect 22560 49292 22612 49298
rect 22560 49234 22612 49240
rect 21640 49224 21692 49230
rect 21640 49166 21692 49172
rect 21824 49224 21876 49230
rect 21824 49166 21876 49172
rect 21088 49088 21140 49094
rect 21088 49030 21140 49036
rect 20628 48204 20680 48210
rect 20628 48146 20680 48152
rect 20996 47660 21048 47666
rect 20996 47602 21048 47608
rect 20272 47110 20392 47138
rect 20456 47518 20576 47546
rect 20272 40769 20300 47110
rect 20352 47048 20404 47054
rect 20352 46990 20404 46996
rect 20364 44266 20392 46990
rect 20352 44260 20404 44266
rect 20352 44202 20404 44208
rect 20258 40760 20314 40769
rect 20258 40695 20314 40704
rect 20456 40610 20484 47518
rect 21008 47462 21036 47602
rect 20536 47456 20588 47462
rect 20536 47398 20588 47404
rect 20996 47456 21048 47462
rect 20996 47398 21048 47404
rect 20548 47122 20576 47398
rect 20536 47116 20588 47122
rect 20536 47058 20588 47064
rect 20536 44260 20588 44266
rect 20536 44202 20588 44208
rect 20272 40582 20484 40610
rect 20166 33008 20222 33017
rect 20166 32943 20222 32952
rect 20168 32836 20220 32842
rect 20168 32778 20220 32784
rect 20180 31210 20208 32778
rect 20272 31890 20300 40582
rect 20444 40520 20496 40526
rect 20350 40488 20406 40497
rect 20444 40462 20496 40468
rect 20350 40423 20406 40432
rect 20260 31884 20312 31890
rect 20260 31826 20312 31832
rect 20260 31408 20312 31414
rect 20260 31350 20312 31356
rect 20168 31204 20220 31210
rect 20168 31146 20220 31152
rect 20180 30802 20208 31146
rect 20272 30841 20300 31350
rect 20258 30832 20314 30841
rect 20168 30796 20220 30802
rect 20258 30767 20314 30776
rect 20168 30738 20220 30744
rect 20168 30660 20220 30666
rect 20168 30602 20220 30608
rect 20076 28756 20128 28762
rect 20076 28698 20128 28704
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 19505 28376 19564 28404
rect 19505 28200 19533 28376
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19984 28212 20036 28218
rect 19505 28172 19564 28200
rect 19432 27872 19484 27878
rect 19432 27814 19484 27820
rect 19536 27554 19564 28172
rect 19984 28154 20036 28160
rect 19708 27872 19760 27878
rect 19708 27814 19760 27820
rect 19444 27526 19564 27554
rect 19340 27396 19392 27402
rect 19340 27338 19392 27344
rect 19352 27130 19380 27338
rect 19340 27124 19392 27130
rect 19340 27066 19392 27072
rect 19444 26858 19472 27526
rect 19720 27470 19748 27814
rect 19708 27464 19760 27470
rect 19706 27432 19708 27441
rect 19760 27432 19762 27441
rect 19996 27402 20024 28154
rect 20088 27674 20116 28426
rect 20076 27668 20128 27674
rect 20076 27610 20128 27616
rect 20074 27432 20130 27441
rect 19706 27367 19762 27376
rect 19984 27396 20036 27402
rect 20074 27367 20130 27376
rect 19984 27338 20036 27344
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19432 26852 19484 26858
rect 19432 26794 19484 26800
rect 19432 26376 19484 26382
rect 19432 26318 19484 26324
rect 19248 26240 19300 26246
rect 19248 26182 19300 26188
rect 19260 25770 19288 26182
rect 19444 25922 19472 26318
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19352 25894 19656 25922
rect 19248 25764 19300 25770
rect 19248 25706 19300 25712
rect 19156 25288 19208 25294
rect 19352 25242 19380 25894
rect 19524 25832 19576 25838
rect 19524 25774 19576 25780
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19444 25362 19472 25638
rect 19432 25356 19484 25362
rect 19432 25298 19484 25304
rect 19536 25294 19564 25774
rect 19628 25702 19656 25894
rect 19616 25696 19668 25702
rect 19616 25638 19668 25644
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19720 25498 19748 25638
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 20088 25362 20116 27367
rect 20076 25356 20128 25362
rect 20076 25298 20128 25304
rect 19156 25230 19208 25236
rect 19168 25158 19196 25230
rect 19260 25214 19380 25242
rect 19524 25288 19576 25294
rect 19524 25230 19576 25236
rect 19156 25152 19208 25158
rect 19156 25094 19208 25100
rect 19260 24834 19288 25214
rect 19340 25152 19392 25158
rect 19340 25094 19392 25100
rect 19984 25152 20036 25158
rect 19984 25094 20036 25100
rect 19168 24818 19288 24834
rect 19352 24818 19380 25094
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 19996 24886 20024 25094
rect 20074 24984 20130 24993
rect 20074 24919 20130 24928
rect 19984 24880 20036 24886
rect 19984 24822 20036 24828
rect 19156 24812 19288 24818
rect 19208 24806 19288 24812
rect 19340 24812 19392 24818
rect 19156 24754 19208 24760
rect 19340 24754 19392 24760
rect 19892 24812 19944 24818
rect 19892 24754 19944 24760
rect 19904 24313 19932 24754
rect 20088 24750 20116 24919
rect 20076 24744 20128 24750
rect 19982 24712 20038 24721
rect 20076 24686 20128 24692
rect 19982 24647 20038 24656
rect 19890 24304 19946 24313
rect 19432 24268 19484 24274
rect 19890 24239 19946 24248
rect 19432 24210 19484 24216
rect 19444 23798 19472 24210
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19156 23792 19208 23798
rect 19156 23734 19208 23740
rect 19432 23792 19484 23798
rect 19432 23734 19484 23740
rect 19168 23118 19196 23734
rect 19444 23526 19472 23734
rect 19432 23520 19484 23526
rect 19432 23462 19484 23468
rect 19156 23112 19208 23118
rect 19156 23054 19208 23060
rect 19168 22642 19196 23054
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19248 22568 19300 22574
rect 19248 22510 19300 22516
rect 19260 21554 19288 22510
rect 19574 21788 19882 21808
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19248 21412 19300 21418
rect 19248 21354 19300 21360
rect 19260 20398 19288 21354
rect 19444 21350 19472 21490
rect 19432 21344 19484 21350
rect 19432 21286 19484 21292
rect 19248 20392 19300 20398
rect 19248 20334 19300 20340
rect 19248 19848 19300 19854
rect 19248 19790 19300 19796
rect 19062 19544 19118 19553
rect 19062 19479 19118 19488
rect 19076 19446 19104 19479
rect 19064 19440 19116 19446
rect 19064 19382 19116 19388
rect 19260 17746 19288 19790
rect 19444 19378 19472 21286
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19892 20256 19944 20262
rect 19892 20198 19944 20204
rect 19904 19854 19932 20198
rect 19892 19848 19944 19854
rect 19892 19790 19944 19796
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19444 18358 19472 19314
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19432 18352 19484 18358
rect 19432 18294 19484 18300
rect 19340 18148 19392 18154
rect 19340 18090 19392 18096
rect 19248 17740 19300 17746
rect 19248 17682 19300 17688
rect 19260 17338 19288 17682
rect 19248 17332 19300 17338
rect 19248 17274 19300 17280
rect 19260 16114 19288 17274
rect 19352 16794 19380 18090
rect 19444 17218 19472 18294
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19444 17190 19564 17218
rect 19432 17060 19484 17066
rect 19432 17002 19484 17008
rect 19340 16788 19392 16794
rect 19340 16730 19392 16736
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19248 16108 19300 16114
rect 19248 16050 19300 16056
rect 19260 15570 19288 16050
rect 19248 15564 19300 15570
rect 19248 15506 19300 15512
rect 19260 13394 19288 15506
rect 19352 14618 19380 16594
rect 19444 16522 19472 17002
rect 19536 16522 19564 17190
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19628 16658 19656 17138
rect 19616 16652 19668 16658
rect 19616 16594 19668 16600
rect 19432 16516 19484 16522
rect 19432 16458 19484 16464
rect 19524 16516 19576 16522
rect 19524 16458 19576 16464
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19444 14958 19472 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19340 14612 19392 14618
rect 19340 14554 19392 14560
rect 19248 13388 19300 13394
rect 19248 13330 19300 13336
rect 19156 13184 19208 13190
rect 19156 13126 19208 13132
rect 19064 11552 19116 11558
rect 19064 11494 19116 11500
rect 19076 11150 19104 11494
rect 19064 11144 19116 11150
rect 19064 11086 19116 11092
rect 19168 10674 19196 13126
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 19260 11150 19288 12786
rect 19352 12238 19380 14554
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19432 13864 19484 13870
rect 19432 13806 19484 13812
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19444 11778 19472 13806
rect 19524 13728 19576 13734
rect 19524 13670 19576 13676
rect 19536 13326 19564 13670
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19444 11750 19564 11778
rect 19248 11144 19300 11150
rect 19248 11086 19300 11092
rect 19156 10668 19208 10674
rect 19156 10610 19208 10616
rect 19064 10464 19116 10470
rect 19064 10406 19116 10412
rect 19076 9586 19104 10406
rect 19260 10062 19288 11086
rect 19536 11082 19564 11750
rect 19616 11756 19668 11762
rect 19616 11698 19668 11704
rect 19628 11354 19656 11698
rect 19616 11348 19668 11354
rect 19616 11290 19668 11296
rect 19996 11234 20024 24647
rect 20074 24440 20130 24449
rect 20074 24375 20130 24384
rect 20088 23730 20116 24375
rect 20076 23724 20128 23730
rect 20076 23666 20128 23672
rect 20076 21548 20128 21554
rect 20076 21490 20128 21496
rect 20088 20466 20116 21490
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20088 19446 20116 20402
rect 20076 19440 20128 19446
rect 20076 19382 20128 19388
rect 20076 17536 20128 17542
rect 20180 17513 20208 30602
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20272 22094 20300 27066
rect 20364 24857 20392 40423
rect 20456 40186 20484 40462
rect 20444 40180 20496 40186
rect 20444 40122 20496 40128
rect 20442 38856 20498 38865
rect 20442 38791 20498 38800
rect 20456 37262 20484 38791
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20444 36304 20496 36310
rect 20444 36246 20496 36252
rect 20456 33386 20484 36246
rect 20444 33380 20496 33386
rect 20444 33322 20496 33328
rect 20444 32904 20496 32910
rect 20444 32846 20496 32852
rect 20456 30870 20484 32846
rect 20444 30864 20496 30870
rect 20444 30806 20496 30812
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20456 26994 20484 27814
rect 20444 26988 20496 26994
rect 20444 26930 20496 26936
rect 20456 26790 20484 26930
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20444 26240 20496 26246
rect 20444 26182 20496 26188
rect 20456 25770 20484 26182
rect 20444 25764 20496 25770
rect 20444 25706 20496 25712
rect 20350 24848 20406 24857
rect 20350 24783 20406 24792
rect 20352 24676 20404 24682
rect 20352 24618 20404 24624
rect 20364 24585 20392 24618
rect 20350 24576 20406 24585
rect 20350 24511 20406 24520
rect 20352 24132 20404 24138
rect 20352 24074 20404 24080
rect 20364 23866 20392 24074
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20352 23656 20404 23662
rect 20350 23624 20352 23633
rect 20404 23624 20406 23633
rect 20350 23559 20406 23568
rect 20272 22066 20392 22094
rect 20258 21992 20314 22001
rect 20258 21927 20260 21936
rect 20312 21927 20314 21936
rect 20260 21898 20312 21904
rect 20260 20528 20312 20534
rect 20260 20470 20312 20476
rect 20272 19990 20300 20470
rect 20260 19984 20312 19990
rect 20260 19926 20312 19932
rect 20260 19848 20312 19854
rect 20260 19790 20312 19796
rect 20076 17478 20128 17484
rect 20166 17504 20222 17513
rect 20088 16726 20116 17478
rect 20166 17439 20222 17448
rect 20076 16720 20128 16726
rect 20272 16674 20300 19790
rect 20364 17542 20392 22066
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20350 17368 20406 17377
rect 20350 17303 20406 17312
rect 20076 16662 20128 16668
rect 20180 16646 20300 16674
rect 20180 14074 20208 16646
rect 20260 16584 20312 16590
rect 20260 16526 20312 16532
rect 20272 14618 20300 16526
rect 20260 14612 20312 14618
rect 20260 14554 20312 14560
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13252 20220 13258
rect 20168 13194 20220 13200
rect 20180 12714 20208 13194
rect 20272 13190 20300 13806
rect 20260 13184 20312 13190
rect 20260 13126 20312 13132
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20168 12708 20220 12714
rect 20168 12650 20220 12656
rect 20168 12164 20220 12170
rect 20168 12106 20220 12112
rect 20180 11898 20208 12106
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20168 11756 20220 11762
rect 20168 11698 20220 11704
rect 20180 11626 20208 11698
rect 20272 11694 20300 12718
rect 20260 11688 20312 11694
rect 20260 11630 20312 11636
rect 20168 11620 20220 11626
rect 20168 11562 20220 11568
rect 19996 11206 20208 11234
rect 19524 11076 19576 11082
rect 19524 11018 19576 11024
rect 19984 11008 20036 11014
rect 20180 10962 20208 11206
rect 19984 10950 20036 10956
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19616 10668 19668 10674
rect 19616 10610 19668 10616
rect 19628 10266 19656 10610
rect 19616 10260 19668 10266
rect 19616 10202 19668 10208
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9586 19288 9998
rect 19340 9988 19392 9994
rect 19340 9930 19392 9936
rect 19064 9580 19116 9586
rect 19064 9522 19116 9528
rect 19248 9580 19300 9586
rect 19248 9522 19300 9528
rect 19260 7970 19288 9522
rect 19352 9382 19380 9930
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19352 8566 19380 9318
rect 19996 9110 20024 10950
rect 20088 10934 20208 10962
rect 19984 9104 20036 9110
rect 19984 9046 20036 9052
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19340 8560 19392 8566
rect 19340 8502 19392 8508
rect 19432 8424 19484 8430
rect 19432 8366 19484 8372
rect 19260 7942 19380 7970
rect 19352 7818 19380 7942
rect 19248 7812 19300 7818
rect 19248 7754 19300 7760
rect 19340 7812 19392 7818
rect 19340 7754 19392 7760
rect 18972 7744 19024 7750
rect 18972 7686 19024 7692
rect 19260 7478 19288 7754
rect 19248 7472 19300 7478
rect 19248 7414 19300 7420
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18696 7268 18748 7274
rect 18696 7210 18748 7216
rect 18328 3596 18380 3602
rect 18328 3538 18380 3544
rect 18144 2848 18196 2854
rect 18144 2790 18196 2796
rect 18708 800 18736 7210
rect 19260 6798 19288 7414
rect 19340 7336 19392 7342
rect 19340 7278 19392 7284
rect 19352 6866 19380 7278
rect 19340 6860 19392 6866
rect 19340 6802 19392 6808
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19444 3738 19472 8366
rect 19996 8090 20024 8910
rect 19984 8084 20036 8090
rect 19984 8026 20036 8032
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 20088 2774 20116 10934
rect 20272 10742 20300 11630
rect 20260 10736 20312 10742
rect 20260 10678 20312 10684
rect 20272 10130 20300 10678
rect 20260 10124 20312 10130
rect 20260 10066 20312 10072
rect 20272 9178 20300 10066
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20180 8362 20208 8910
rect 20168 8356 20220 8362
rect 20168 8298 20220 8304
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20272 3058 20300 3470
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20088 2746 20208 2774
rect 20180 2582 20208 2746
rect 20364 2582 20392 17303
rect 20456 11898 20484 25706
rect 20548 22094 20576 44202
rect 20720 42152 20772 42158
rect 20720 42094 20772 42100
rect 20732 41002 20760 42094
rect 20904 41472 20956 41478
rect 20904 41414 20956 41420
rect 20916 41138 20944 41414
rect 20904 41132 20956 41138
rect 20904 41074 20956 41080
rect 20812 41064 20864 41070
rect 20812 41006 20864 41012
rect 20720 40996 20772 41002
rect 20720 40938 20772 40944
rect 20824 40390 20852 41006
rect 20812 40384 20864 40390
rect 20812 40326 20864 40332
rect 20628 39908 20680 39914
rect 20628 39850 20680 39856
rect 20640 37262 20668 39850
rect 20824 39506 20852 40326
rect 20812 39500 20864 39506
rect 20812 39442 20864 39448
rect 20720 39432 20772 39438
rect 20718 39400 20720 39409
rect 20772 39400 20774 39409
rect 20718 39335 20774 39344
rect 20732 39098 20760 39335
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 20916 38865 20944 41074
rect 20902 38856 20958 38865
rect 20902 38791 20958 38800
rect 21100 38350 21128 49030
rect 21836 48754 21864 49166
rect 22284 49156 22336 49162
rect 22284 49098 22336 49104
rect 21824 48748 21876 48754
rect 21824 48690 21876 48696
rect 22296 47802 22324 49098
rect 22376 49088 22428 49094
rect 23400 49076 23428 51326
rect 23846 51200 23902 52000
rect 24490 51200 24546 52000
rect 25134 51200 25190 52000
rect 25778 51354 25834 52000
rect 25778 51326 26004 51354
rect 25778 51200 25834 51326
rect 23860 49230 23888 51200
rect 24124 49360 24176 49366
rect 24124 49302 24176 49308
rect 23848 49224 23900 49230
rect 23848 49166 23900 49172
rect 23400 49048 23520 49076
rect 22376 49030 22428 49036
rect 22284 47796 22336 47802
rect 22284 47738 22336 47744
rect 21364 45824 21416 45830
rect 21364 45766 21416 45772
rect 21272 38548 21324 38554
rect 21272 38490 21324 38496
rect 21088 38344 21140 38350
rect 21088 38286 21140 38292
rect 21180 37800 21232 37806
rect 21180 37742 21232 37748
rect 20996 37732 21048 37738
rect 20996 37674 21048 37680
rect 20628 37256 20680 37262
rect 20628 37198 20680 37204
rect 20640 36650 20668 37198
rect 21008 36718 21036 37674
rect 21088 37664 21140 37670
rect 21088 37606 21140 37612
rect 21100 37262 21128 37606
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 21192 36922 21220 37742
rect 21180 36916 21232 36922
rect 21180 36858 21232 36864
rect 20996 36712 21048 36718
rect 20996 36654 21048 36660
rect 20628 36644 20680 36650
rect 20628 36586 20680 36592
rect 20640 32502 20668 36586
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 20916 36242 20944 36518
rect 20904 36236 20956 36242
rect 20904 36178 20956 36184
rect 20720 35760 20772 35766
rect 20718 35728 20720 35737
rect 20772 35728 20774 35737
rect 21008 35698 21036 36654
rect 21088 36032 21140 36038
rect 21088 35974 21140 35980
rect 21100 35698 21128 35974
rect 20718 35663 20774 35672
rect 20812 35692 20864 35698
rect 20996 35692 21048 35698
rect 20864 35652 20944 35680
rect 20812 35634 20864 35640
rect 20720 35012 20772 35018
rect 20720 34954 20772 34960
rect 20732 34746 20760 34954
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20812 32972 20864 32978
rect 20812 32914 20864 32920
rect 20720 32768 20772 32774
rect 20720 32710 20772 32716
rect 20628 32496 20680 32502
rect 20628 32438 20680 32444
rect 20628 31408 20680 31414
rect 20732 31396 20760 32710
rect 20680 31368 20760 31396
rect 20628 31350 20680 31356
rect 20824 31278 20852 32914
rect 20812 31272 20864 31278
rect 20812 31214 20864 31220
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20824 29646 20852 30534
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20628 29572 20680 29578
rect 20628 29514 20680 29520
rect 20640 26382 20668 29514
rect 20812 28416 20864 28422
rect 20810 28384 20812 28393
rect 20864 28384 20866 28393
rect 20810 28319 20866 28328
rect 20824 27062 20852 28319
rect 20812 27056 20864 27062
rect 20812 26998 20864 27004
rect 20628 26376 20680 26382
rect 20628 26318 20680 26324
rect 20812 25220 20864 25226
rect 20812 25162 20864 25168
rect 20824 24936 20852 25162
rect 20640 24908 20852 24936
rect 20640 24682 20668 24908
rect 20803 24812 20855 24818
rect 20732 24772 20803 24800
rect 20628 24676 20680 24682
rect 20628 24618 20680 24624
rect 20732 24562 20760 24772
rect 20803 24754 20855 24760
rect 20640 24534 20760 24562
rect 20640 24070 20668 24534
rect 20628 24064 20680 24070
rect 20628 24006 20680 24012
rect 20720 24064 20772 24070
rect 20720 24006 20772 24012
rect 20640 23594 20668 24006
rect 20628 23588 20680 23594
rect 20628 23530 20680 23536
rect 20732 23050 20760 24006
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20824 23254 20852 23666
rect 20812 23248 20864 23254
rect 20812 23190 20864 23196
rect 20720 23044 20772 23050
rect 20720 22986 20772 22992
rect 20812 23044 20864 23050
rect 20812 22986 20864 22992
rect 20720 22228 20772 22234
rect 20720 22170 20772 22176
rect 20548 22066 20668 22094
rect 20640 21978 20668 22066
rect 20732 22030 20760 22170
rect 20548 21950 20668 21978
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20548 19990 20576 21950
rect 20628 21888 20680 21894
rect 20628 21830 20680 21836
rect 20640 21622 20668 21830
rect 20824 21622 20852 22986
rect 20628 21616 20680 21622
rect 20812 21616 20864 21622
rect 20628 21558 20680 21564
rect 20718 21584 20774 21593
rect 20812 21558 20864 21564
rect 20718 21519 20774 21528
rect 20732 20942 20760 21519
rect 20720 20936 20772 20942
rect 20720 20878 20772 20884
rect 20732 20618 20760 20878
rect 20732 20590 20852 20618
rect 20720 20460 20772 20466
rect 20720 20402 20772 20408
rect 20536 19984 20588 19990
rect 20536 19926 20588 19932
rect 20732 19242 20760 20402
rect 20720 19236 20772 19242
rect 20720 19178 20772 19184
rect 20536 19168 20588 19174
rect 20536 19110 20588 19116
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20444 11076 20496 11082
rect 20444 11018 20496 11024
rect 20456 2922 20484 11018
rect 20444 2916 20496 2922
rect 20444 2858 20496 2864
rect 20168 2576 20220 2582
rect 20168 2518 20220 2524
rect 20352 2576 20404 2582
rect 20352 2518 20404 2524
rect 20548 2446 20576 19110
rect 20626 18320 20682 18329
rect 20626 18255 20628 18264
rect 20680 18255 20682 18264
rect 20628 18226 20680 18232
rect 20640 17882 20668 18226
rect 20628 17876 20680 17882
rect 20628 17818 20680 17824
rect 20824 17678 20852 20590
rect 20812 17672 20864 17678
rect 20812 17614 20864 17620
rect 20628 17604 20680 17610
rect 20628 17546 20680 17552
rect 20640 16998 20668 17546
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20628 16584 20680 16590
rect 20628 16526 20680 16532
rect 20640 15978 20668 16526
rect 20628 15972 20680 15978
rect 20628 15914 20680 15920
rect 20824 14414 20852 17614
rect 20812 14408 20864 14414
rect 20812 14350 20864 14356
rect 20824 14090 20852 14350
rect 20732 14062 20852 14090
rect 20732 13938 20760 14062
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 11892 20680 11898
rect 20628 11834 20680 11840
rect 20640 10674 20668 11834
rect 20732 11762 20760 12582
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20720 11756 20772 11762
rect 20720 11698 20772 11704
rect 20628 10668 20680 10674
rect 20628 10610 20680 10616
rect 20640 10198 20668 10610
rect 20628 10192 20680 10198
rect 20628 10134 20680 10140
rect 20720 10056 20772 10062
rect 20720 9998 20772 10004
rect 20824 10010 20852 11834
rect 20916 11506 20944 35652
rect 20996 35634 21048 35640
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21008 35018 21036 35634
rect 21284 35154 21312 38490
rect 21272 35148 21324 35154
rect 21272 35090 21324 35096
rect 20996 35012 21048 35018
rect 20996 34954 21048 34960
rect 21272 34536 21324 34542
rect 21272 34478 21324 34484
rect 21284 34066 21312 34478
rect 21272 34060 21324 34066
rect 21272 34002 21324 34008
rect 21284 33590 21312 34002
rect 21272 33584 21324 33590
rect 21272 33526 21324 33532
rect 21088 32768 21140 32774
rect 21088 32710 21140 32716
rect 21100 32570 21128 32710
rect 21088 32564 21140 32570
rect 21088 32506 21140 32512
rect 21088 31884 21140 31890
rect 21088 31826 21140 31832
rect 20996 31816 21048 31822
rect 20996 31758 21048 31764
rect 21008 31482 21036 31758
rect 20996 31476 21048 31482
rect 20996 31418 21048 31424
rect 21008 31346 21036 31418
rect 20996 31340 21048 31346
rect 20996 31282 21048 31288
rect 21008 30258 21036 31282
rect 21100 30297 21128 31826
rect 21376 31754 21404 45766
rect 22388 44690 22416 49030
rect 23492 48686 23520 49048
rect 22652 48680 22704 48686
rect 22652 48622 22704 48628
rect 23480 48680 23532 48686
rect 23480 48622 23532 48628
rect 22664 48346 22692 48622
rect 22652 48340 22704 48346
rect 22652 48282 22704 48288
rect 23664 48136 23716 48142
rect 23664 48078 23716 48084
rect 23572 48068 23624 48074
rect 23572 48010 23624 48016
rect 23584 47734 23612 48010
rect 23572 47728 23624 47734
rect 23572 47670 23624 47676
rect 22560 47660 22612 47666
rect 22560 47602 22612 47608
rect 22296 44662 22416 44690
rect 21916 43852 21968 43858
rect 21916 43794 21968 43800
rect 21824 41540 21876 41546
rect 21824 41482 21876 41488
rect 21836 41274 21864 41482
rect 21824 41268 21876 41274
rect 21824 41210 21876 41216
rect 21928 41206 21956 43794
rect 22192 41472 22244 41478
rect 22192 41414 22244 41420
rect 21916 41200 21968 41206
rect 21916 41142 21968 41148
rect 22204 40610 22232 41414
rect 22296 41274 22324 44662
rect 22376 41540 22428 41546
rect 22376 41482 22428 41488
rect 22284 41268 22336 41274
rect 22284 41210 22336 41216
rect 22284 41132 22336 41138
rect 22284 41074 22336 41080
rect 22296 40730 22324 41074
rect 22388 41070 22416 41482
rect 22376 41064 22428 41070
rect 22376 41006 22428 41012
rect 22284 40724 22336 40730
rect 22284 40666 22336 40672
rect 22112 40582 22232 40610
rect 22112 40526 22140 40582
rect 22100 40520 22152 40526
rect 22100 40462 22152 40468
rect 22112 38418 22140 40462
rect 22192 39976 22244 39982
rect 22192 39918 22244 39924
rect 22100 38412 22152 38418
rect 22100 38354 22152 38360
rect 22008 38208 22060 38214
rect 22008 38150 22060 38156
rect 22020 37942 22048 38150
rect 22008 37936 22060 37942
rect 22008 37878 22060 37884
rect 22204 37806 22232 39918
rect 22284 38888 22336 38894
rect 22282 38856 22284 38865
rect 22336 38856 22338 38865
rect 22282 38791 22338 38800
rect 22376 38344 22428 38350
rect 22428 38304 22508 38332
rect 22376 38286 22428 38292
rect 22376 37868 22428 37874
rect 22376 37810 22428 37816
rect 22192 37800 22244 37806
rect 22192 37742 22244 37748
rect 22204 36378 22232 37742
rect 22192 36372 22244 36378
rect 22192 36314 22244 36320
rect 22204 35766 22232 36314
rect 22388 36145 22416 37810
rect 22480 36310 22508 38304
rect 22468 36304 22520 36310
rect 22468 36246 22520 36252
rect 22374 36136 22430 36145
rect 22374 36071 22430 36080
rect 22192 35760 22244 35766
rect 21914 35728 21970 35737
rect 21456 35692 21508 35698
rect 22192 35702 22244 35708
rect 21914 35663 21916 35672
rect 21456 35634 21508 35640
rect 21968 35663 21970 35672
rect 21916 35634 21968 35640
rect 21468 35057 21496 35634
rect 22006 35456 22062 35465
rect 22006 35391 22062 35400
rect 22020 35086 22048 35391
rect 21548 35080 21600 35086
rect 21454 35048 21510 35057
rect 21916 35080 21968 35086
rect 21600 35040 21680 35068
rect 21548 35022 21600 35028
rect 21454 34983 21510 34992
rect 21652 32042 21680 35040
rect 21914 35048 21916 35057
rect 22008 35080 22060 35086
rect 21968 35048 21970 35057
rect 21836 35006 21914 35034
rect 21836 33998 21864 35006
rect 22008 35022 22060 35028
rect 21914 34983 21970 34992
rect 21916 34944 21968 34950
rect 21916 34886 21968 34892
rect 21928 34610 21956 34886
rect 21916 34604 21968 34610
rect 21916 34546 21968 34552
rect 21824 33992 21876 33998
rect 21824 33934 21876 33940
rect 21824 32972 21876 32978
rect 21824 32914 21876 32920
rect 21652 32014 21772 32042
rect 21376 31726 21588 31754
rect 21364 31204 21416 31210
rect 21364 31146 21416 31152
rect 21376 30666 21404 31146
rect 21272 30660 21324 30666
rect 21272 30602 21324 30608
rect 21364 30660 21416 30666
rect 21364 30602 21416 30608
rect 21284 30394 21312 30602
rect 21272 30388 21324 30394
rect 21272 30330 21324 30336
rect 21086 30288 21142 30297
rect 20996 30252 21048 30258
rect 21086 30223 21142 30232
rect 20996 30194 21048 30200
rect 21088 29164 21140 29170
rect 21088 29106 21140 29112
rect 20996 28756 21048 28762
rect 20996 28698 21048 28704
rect 21008 27418 21036 28698
rect 21100 27606 21128 29106
rect 21088 27600 21140 27606
rect 21088 27542 21140 27548
rect 21008 27390 21128 27418
rect 20996 24744 21048 24750
rect 20996 24686 21048 24692
rect 21008 23866 21036 24686
rect 20996 23860 21048 23866
rect 20996 23802 21048 23808
rect 20996 22024 21048 22030
rect 20996 21966 21048 21972
rect 21008 21729 21036 21966
rect 20994 21720 21050 21729
rect 20994 21655 21050 21664
rect 20996 21616 21048 21622
rect 20996 21558 21048 21564
rect 21008 21146 21036 21558
rect 20996 21140 21048 21146
rect 20996 21082 21048 21088
rect 20996 20800 21048 20806
rect 20996 20742 21048 20748
rect 21008 20466 21036 20742
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20996 15360 21048 15366
rect 20996 15302 21048 15308
rect 21008 14958 21036 15302
rect 20996 14952 21048 14958
rect 20996 14894 21048 14900
rect 21008 13870 21036 14894
rect 20996 13864 21048 13870
rect 20996 13806 21048 13812
rect 21100 11898 21128 27390
rect 21272 27396 21324 27402
rect 21272 27338 21324 27344
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21192 24449 21220 24754
rect 21178 24440 21234 24449
rect 21178 24375 21234 24384
rect 21192 23730 21220 24375
rect 21180 23724 21232 23730
rect 21180 23666 21232 23672
rect 21180 22976 21232 22982
rect 21180 22918 21232 22924
rect 21192 22710 21220 22918
rect 21180 22704 21232 22710
rect 21180 22646 21232 22652
rect 21192 21593 21220 22646
rect 21178 21584 21234 21593
rect 21178 21519 21234 21528
rect 21180 21480 21232 21486
rect 21180 21422 21232 21428
rect 21192 19854 21220 21422
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21192 19310 21220 19790
rect 21180 19304 21232 19310
rect 21180 19246 21232 19252
rect 21192 18290 21220 19246
rect 21180 18284 21232 18290
rect 21180 18226 21232 18232
rect 21284 16590 21312 27338
rect 21560 25362 21588 31726
rect 21640 30592 21692 30598
rect 21640 30534 21692 30540
rect 21652 30326 21680 30534
rect 21640 30320 21692 30326
rect 21640 30262 21692 30268
rect 21548 25356 21600 25362
rect 21548 25298 21600 25304
rect 21548 25152 21600 25158
rect 21548 25094 21600 25100
rect 21364 24812 21416 24818
rect 21364 24754 21416 24760
rect 21376 24721 21404 24754
rect 21362 24712 21418 24721
rect 21362 24647 21418 24656
rect 21560 23526 21588 25094
rect 21640 24676 21692 24682
rect 21640 24618 21692 24624
rect 21652 24585 21680 24618
rect 21638 24576 21694 24585
rect 21638 24511 21694 24520
rect 21744 24290 21772 32014
rect 21836 30802 21864 32914
rect 22020 32842 22048 35022
rect 22204 34678 22232 35702
rect 22192 34672 22244 34678
rect 22192 34614 22244 34620
rect 22284 33924 22336 33930
rect 22284 33866 22336 33872
rect 22296 33590 22324 33866
rect 22388 33658 22416 36071
rect 22376 33652 22428 33658
rect 22376 33594 22428 33600
rect 22284 33584 22336 33590
rect 22388 33561 22416 33594
rect 22284 33526 22336 33532
rect 22374 33552 22430 33561
rect 22100 33448 22152 33454
rect 22100 33390 22152 33396
rect 22008 32836 22060 32842
rect 22008 32778 22060 32784
rect 21916 32428 21968 32434
rect 21916 32370 21968 32376
rect 21928 32026 21956 32370
rect 21916 32020 21968 32026
rect 21916 31962 21968 31968
rect 22008 31748 22060 31754
rect 22112 31736 22140 33390
rect 22192 32768 22244 32774
rect 22192 32710 22244 32716
rect 22060 31708 22140 31736
rect 22008 31690 22060 31696
rect 22204 31414 22232 32710
rect 22296 32502 22324 33526
rect 22374 33487 22430 33496
rect 22480 33454 22508 36246
rect 22468 33448 22520 33454
rect 22468 33390 22520 33396
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22388 31482 22416 31758
rect 22468 31680 22520 31686
rect 22468 31622 22520 31628
rect 22480 31482 22508 31622
rect 22376 31476 22428 31482
rect 22376 31418 22428 31424
rect 22468 31476 22520 31482
rect 22468 31418 22520 31424
rect 22192 31408 22244 31414
rect 22192 31350 22244 31356
rect 21824 30796 21876 30802
rect 22572 30784 22600 47602
rect 23676 46646 23704 48078
rect 24032 48000 24084 48006
rect 24032 47942 24084 47948
rect 24044 47258 24072 47942
rect 24032 47252 24084 47258
rect 24032 47194 24084 47200
rect 23664 46640 23716 46646
rect 23664 46582 23716 46588
rect 23388 43444 23440 43450
rect 23388 43386 23440 43392
rect 22928 42220 22980 42226
rect 22928 42162 22980 42168
rect 22652 40588 22704 40594
rect 22652 40530 22704 40536
rect 22664 39982 22692 40530
rect 22940 40526 22968 42162
rect 23020 41540 23072 41546
rect 23020 41482 23072 41488
rect 22928 40520 22980 40526
rect 22928 40462 22980 40468
rect 22940 40390 22968 40462
rect 22928 40384 22980 40390
rect 22928 40326 22980 40332
rect 22928 40180 22980 40186
rect 22928 40122 22980 40128
rect 22836 40044 22888 40050
rect 22836 39986 22888 39992
rect 22652 39976 22704 39982
rect 22652 39918 22704 39924
rect 22848 39642 22876 39986
rect 22836 39636 22888 39642
rect 22836 39578 22888 39584
rect 22940 38554 22968 40122
rect 23032 39302 23060 41482
rect 23204 41064 23256 41070
rect 23204 41006 23256 41012
rect 23216 40594 23244 41006
rect 23204 40588 23256 40594
rect 23204 40530 23256 40536
rect 23112 40452 23164 40458
rect 23112 40394 23164 40400
rect 23124 39438 23152 40394
rect 23112 39432 23164 39438
rect 23112 39374 23164 39380
rect 23020 39296 23072 39302
rect 23020 39238 23072 39244
rect 22928 38548 22980 38554
rect 22928 38490 22980 38496
rect 23112 38412 23164 38418
rect 23112 38354 23164 38360
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 37942 22876 38286
rect 23020 38276 23072 38282
rect 23020 38218 23072 38224
rect 22836 37936 22888 37942
rect 22836 37878 22888 37884
rect 23032 37466 23060 38218
rect 23020 37460 23072 37466
rect 23020 37402 23072 37408
rect 22744 37324 22796 37330
rect 22744 37266 22796 37272
rect 22756 37126 22784 37266
rect 22744 37120 22796 37126
rect 22744 37062 22796 37068
rect 22756 34202 22784 37062
rect 23124 36174 23152 38354
rect 23112 36168 23164 36174
rect 23112 36110 23164 36116
rect 23112 36032 23164 36038
rect 23112 35974 23164 35980
rect 23204 36032 23256 36038
rect 23204 35974 23256 35980
rect 23124 34898 23152 35974
rect 23216 35154 23244 35974
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23308 35154 23336 35430
rect 23204 35148 23256 35154
rect 23204 35090 23256 35096
rect 23296 35148 23348 35154
rect 23296 35090 23348 35096
rect 23308 34898 23336 35090
rect 23124 34870 23336 34898
rect 22836 34740 22888 34746
rect 22836 34682 22888 34688
rect 22744 34196 22796 34202
rect 22744 34138 22796 34144
rect 22652 31884 22704 31890
rect 22652 31826 22704 31832
rect 21824 30738 21876 30744
rect 22388 30756 22600 30784
rect 22100 30728 22152 30734
rect 22100 30670 22152 30676
rect 22112 29492 22140 30670
rect 22192 29504 22244 29510
rect 22112 29464 22192 29492
rect 22192 29446 22244 29452
rect 22204 29306 22232 29446
rect 22192 29300 22244 29306
rect 22192 29242 22244 29248
rect 22284 28484 22336 28490
rect 22284 28426 22336 28432
rect 22192 25220 22244 25226
rect 22192 25162 22244 25168
rect 21744 24262 22048 24290
rect 21824 24200 21876 24206
rect 21824 24142 21876 24148
rect 21640 24132 21692 24138
rect 21640 24074 21692 24080
rect 21732 24132 21784 24138
rect 21732 24074 21784 24080
rect 21548 23520 21600 23526
rect 21548 23462 21600 23468
rect 21364 22500 21416 22506
rect 21364 22442 21416 22448
rect 21376 17218 21404 22442
rect 21548 21548 21600 21554
rect 21548 21490 21600 21496
rect 21560 21078 21588 21490
rect 21548 21072 21600 21078
rect 21548 21014 21600 21020
rect 21456 21004 21508 21010
rect 21456 20946 21508 20952
rect 21468 20806 21496 20946
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21456 20256 21508 20262
rect 21456 20198 21508 20204
rect 21468 19854 21496 20198
rect 21456 19848 21508 19854
rect 21456 19790 21508 19796
rect 21376 17190 21588 17218
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21456 14544 21508 14550
rect 21456 14486 21508 14492
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21088 11892 21140 11898
rect 21088 11834 21140 11840
rect 21192 11608 21220 14214
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21272 12844 21324 12850
rect 21272 12786 21324 12792
rect 21284 12442 21312 12786
rect 21272 12436 21324 12442
rect 21272 12378 21324 12384
rect 21284 11830 21312 12378
rect 21376 12238 21404 13262
rect 21364 12232 21416 12238
rect 21364 12174 21416 12180
rect 21272 11824 21324 11830
rect 21272 11766 21324 11772
rect 21192 11580 21312 11608
rect 20916 11478 21220 11506
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 20732 9722 20760 9998
rect 20824 9982 21036 10010
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20720 9716 20772 9722
rect 20720 9658 20772 9664
rect 20916 8974 20944 9862
rect 20720 8968 20772 8974
rect 20720 8910 20772 8916
rect 20904 8968 20956 8974
rect 20904 8910 20956 8916
rect 20732 8838 20760 8910
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20720 8832 20772 8838
rect 20720 8774 20772 8780
rect 20824 8430 20852 8842
rect 20812 8424 20864 8430
rect 20812 8366 20864 8372
rect 20720 8084 20772 8090
rect 20720 8026 20772 8032
rect 20732 6798 20760 8026
rect 20904 7744 20956 7750
rect 20904 7686 20956 7692
rect 20812 7404 20864 7410
rect 20812 7346 20864 7352
rect 20824 6866 20852 7346
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20916 6798 20944 7686
rect 20720 6792 20772 6798
rect 20720 6734 20772 6740
rect 20904 6792 20956 6798
rect 20904 6734 20956 6740
rect 21008 6746 21036 9982
rect 21100 9654 21128 11086
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21100 8838 21128 9590
rect 21088 8832 21140 8838
rect 21088 8774 21140 8780
rect 21100 7342 21128 8774
rect 21088 7336 21140 7342
rect 21088 7278 21140 7284
rect 21100 6866 21128 7278
rect 21088 6860 21140 6866
rect 21088 6802 21140 6808
rect 21008 6718 21128 6746
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20628 3596 20680 3602
rect 20628 3538 20680 3544
rect 20536 2440 20588 2446
rect 20536 2382 20588 2388
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 19996 800 20024 2314
rect 20640 800 20668 3538
rect 21008 2514 21036 3878
rect 20996 2508 21048 2514
rect 20996 2450 21048 2456
rect 21100 2378 21128 6718
rect 21088 2372 21140 2378
rect 21088 2314 21140 2320
rect 21192 2038 21220 11478
rect 21284 11014 21312 11580
rect 21376 11150 21404 12174
rect 21364 11144 21416 11150
rect 21364 11086 21416 11092
rect 21272 11008 21324 11014
rect 21272 10950 21324 10956
rect 21468 8106 21496 14486
rect 21560 11558 21588 17190
rect 21548 11552 21600 11558
rect 21548 11494 21600 11500
rect 21560 10266 21588 11494
rect 21548 10260 21600 10266
rect 21548 10202 21600 10208
rect 21376 8078 21588 8106
rect 21376 8022 21404 8078
rect 21364 8016 21416 8022
rect 21364 7958 21416 7964
rect 21456 7744 21508 7750
rect 21456 7686 21508 7692
rect 21468 6730 21496 7686
rect 21456 6724 21508 6730
rect 21456 6666 21508 6672
rect 21560 6662 21588 8078
rect 21548 6656 21600 6662
rect 21548 6598 21600 6604
rect 21652 2650 21680 24074
rect 21744 23050 21772 24074
rect 21732 23044 21784 23050
rect 21732 22986 21784 22992
rect 21836 22642 21864 24142
rect 21916 23588 21968 23594
rect 21916 23530 21968 23536
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21732 22432 21784 22438
rect 21732 22374 21784 22380
rect 21744 22030 21772 22374
rect 21836 22234 21864 22578
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21732 22024 21784 22030
rect 21732 21966 21784 21972
rect 21836 21486 21864 22170
rect 21928 22098 21956 23530
rect 21916 22092 21968 22098
rect 21916 22034 21968 22040
rect 21824 21480 21876 21486
rect 21824 21422 21876 21428
rect 21732 20392 21784 20398
rect 21732 20334 21784 20340
rect 21744 14550 21772 20334
rect 21916 20256 21968 20262
rect 21916 20198 21968 20204
rect 21822 17912 21878 17921
rect 21822 17847 21878 17856
rect 21732 14544 21784 14550
rect 21732 14486 21784 14492
rect 21836 13530 21864 17847
rect 21824 13524 21876 13530
rect 21824 13466 21876 13472
rect 21928 12434 21956 20198
rect 21744 12406 21956 12434
rect 21744 8090 21772 12406
rect 21916 11552 21968 11558
rect 21916 11494 21968 11500
rect 21928 11150 21956 11494
rect 21916 11144 21968 11150
rect 21916 11086 21968 11092
rect 21916 9580 21968 9586
rect 21916 9522 21968 9528
rect 21928 8838 21956 9522
rect 21916 8832 21968 8838
rect 21916 8774 21968 8780
rect 21824 8424 21876 8430
rect 21824 8366 21876 8372
rect 21732 8084 21784 8090
rect 21732 8026 21784 8032
rect 21744 7886 21772 8026
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21836 7002 21864 8366
rect 21824 6996 21876 7002
rect 21824 6938 21876 6944
rect 21928 4690 21956 8774
rect 21916 4684 21968 4690
rect 21916 4626 21968 4632
rect 22020 2774 22048 24262
rect 22100 22636 22152 22642
rect 22100 22578 22152 22584
rect 22112 22001 22140 22578
rect 22098 21992 22154 22001
rect 22098 21927 22154 21936
rect 22100 20936 22152 20942
rect 22100 20878 22152 20884
rect 22112 20466 22140 20878
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22204 19174 22232 25162
rect 22296 22166 22324 28426
rect 22388 25770 22416 30756
rect 22560 27600 22612 27606
rect 22560 27542 22612 27548
rect 22572 27418 22600 27542
rect 22480 27390 22600 27418
rect 22480 27334 22508 27390
rect 22468 27328 22520 27334
rect 22468 27270 22520 27276
rect 22560 27328 22612 27334
rect 22560 27270 22612 27276
rect 22572 26994 22600 27270
rect 22560 26988 22612 26994
rect 22560 26930 22612 26936
rect 22376 25764 22428 25770
rect 22376 25706 22428 25712
rect 22284 22160 22336 22166
rect 22284 22102 22336 22108
rect 22664 22094 22692 31826
rect 22756 30598 22784 34138
rect 22744 30592 22796 30598
rect 22744 30534 22796 30540
rect 22744 30048 22796 30054
rect 22744 29990 22796 29996
rect 22756 29782 22784 29990
rect 22744 29776 22796 29782
rect 22744 29718 22796 29724
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22756 27062 22784 27814
rect 22744 27056 22796 27062
rect 22744 26998 22796 27004
rect 22848 24410 22876 34682
rect 22928 32836 22980 32842
rect 22928 32778 22980 32784
rect 22940 32230 22968 32778
rect 23124 32774 23152 34870
rect 23400 32960 23428 43386
rect 23572 42016 23624 42022
rect 23572 41958 23624 41964
rect 23584 41614 23612 41958
rect 23572 41608 23624 41614
rect 23572 41550 23624 41556
rect 23756 41608 23808 41614
rect 23756 41550 23808 41556
rect 23480 41472 23532 41478
rect 23480 41414 23532 41420
rect 23492 41206 23520 41414
rect 23480 41200 23532 41206
rect 23480 41142 23532 41148
rect 23768 41138 23796 41550
rect 23756 41132 23808 41138
rect 23756 41074 23808 41080
rect 23768 40118 23796 41074
rect 23756 40112 23808 40118
rect 23756 40054 23808 40060
rect 23768 39370 23796 40054
rect 24136 40050 24164 49302
rect 24504 48278 24532 51200
rect 25976 49230 26004 51326
rect 26422 51200 26478 52000
rect 27066 51200 27122 52000
rect 27710 51354 27766 52000
rect 28354 51354 28410 52000
rect 27710 51326 27844 51354
rect 27710 51200 27766 51326
rect 26436 49230 26464 51200
rect 25964 49224 26016 49230
rect 25964 49166 26016 49172
rect 26424 49224 26476 49230
rect 26424 49166 26476 49172
rect 25412 49088 25464 49094
rect 25412 49030 25464 49036
rect 24952 48544 25004 48550
rect 24952 48486 25004 48492
rect 24492 48272 24544 48278
rect 24492 48214 24544 48220
rect 24964 48210 24992 48486
rect 24952 48204 25004 48210
rect 24952 48146 25004 48152
rect 24768 46640 24820 46646
rect 24768 46582 24820 46588
rect 24584 42220 24636 42226
rect 24584 42162 24636 42168
rect 24596 41018 24624 42162
rect 24596 40990 24716 41018
rect 24688 40934 24716 40990
rect 24676 40928 24728 40934
rect 24676 40870 24728 40876
rect 24584 40452 24636 40458
rect 24584 40394 24636 40400
rect 24492 40384 24544 40390
rect 24492 40326 24544 40332
rect 24124 40044 24176 40050
rect 24124 39986 24176 39992
rect 23848 39976 23900 39982
rect 23848 39918 23900 39924
rect 23860 39438 23888 39918
rect 24504 39438 24532 40326
rect 24596 40186 24624 40394
rect 24584 40180 24636 40186
rect 24584 40122 24636 40128
rect 23848 39432 23900 39438
rect 23848 39374 23900 39380
rect 24492 39432 24544 39438
rect 24492 39374 24544 39380
rect 23756 39364 23808 39370
rect 23756 39306 23808 39312
rect 23860 39098 23888 39374
rect 24032 39296 24084 39302
rect 24032 39238 24084 39244
rect 23848 39092 23900 39098
rect 23848 39034 23900 39040
rect 24044 39030 24072 39238
rect 24032 39024 24084 39030
rect 24032 38966 24084 38972
rect 24216 38956 24268 38962
rect 24216 38898 24268 38904
rect 24228 38418 24256 38898
rect 24216 38412 24268 38418
rect 24216 38354 24268 38360
rect 23572 38344 23624 38350
rect 23572 38286 23624 38292
rect 23584 36786 23612 38286
rect 23756 37188 23808 37194
rect 23756 37130 23808 37136
rect 23768 36786 23796 37130
rect 23572 36780 23624 36786
rect 23572 36722 23624 36728
rect 23756 36780 23808 36786
rect 23756 36722 23808 36728
rect 23584 36650 23612 36722
rect 23572 36644 23624 36650
rect 23572 36586 23624 36592
rect 23664 35692 23716 35698
rect 23664 35634 23716 35640
rect 23480 35012 23532 35018
rect 23480 34954 23532 34960
rect 23492 34678 23520 34954
rect 23480 34672 23532 34678
rect 23480 34614 23532 34620
rect 23676 34542 23704 35634
rect 23768 35630 23796 36722
rect 24228 35766 24256 38354
rect 24308 37664 24360 37670
rect 24308 37606 24360 37612
rect 24320 37262 24348 37606
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24412 36854 24440 37062
rect 24400 36848 24452 36854
rect 24400 36790 24452 36796
rect 24400 36100 24452 36106
rect 24400 36042 24452 36048
rect 24216 35760 24268 35766
rect 24216 35702 24268 35708
rect 23756 35624 23808 35630
rect 23756 35566 23808 35572
rect 23768 34542 23796 35566
rect 23664 34536 23716 34542
rect 23664 34478 23716 34484
rect 23756 34536 23808 34542
rect 23756 34478 23808 34484
rect 23480 34400 23532 34406
rect 23480 34342 23532 34348
rect 23492 33930 23520 34342
rect 23768 33930 23796 34478
rect 23940 34128 23992 34134
rect 23940 34070 23992 34076
rect 23480 33924 23532 33930
rect 23480 33866 23532 33872
rect 23756 33924 23808 33930
rect 23756 33866 23808 33872
rect 23572 33856 23624 33862
rect 23572 33798 23624 33804
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23584 33658 23612 33798
rect 23572 33652 23624 33658
rect 23572 33594 23624 33600
rect 23860 33522 23888 33798
rect 23572 33516 23624 33522
rect 23848 33516 23900 33522
rect 23624 33476 23704 33504
rect 23572 33458 23624 33464
rect 23480 33380 23532 33386
rect 23480 33322 23532 33328
rect 23216 32932 23428 32960
rect 23112 32768 23164 32774
rect 23112 32710 23164 32716
rect 22928 32224 22980 32230
rect 22928 32166 22980 32172
rect 23020 31340 23072 31346
rect 23020 31282 23072 31288
rect 23032 30938 23060 31282
rect 23112 31272 23164 31278
rect 23112 31214 23164 31220
rect 23020 30932 23072 30938
rect 23020 30874 23072 30880
rect 23124 30734 23152 31214
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 23032 30258 23060 30534
rect 23020 30252 23072 30258
rect 23020 30194 23072 30200
rect 23112 29096 23164 29102
rect 23112 29038 23164 29044
rect 23124 28082 23152 29038
rect 23112 28076 23164 28082
rect 23112 28018 23164 28024
rect 23020 27328 23072 27334
rect 23020 27270 23072 27276
rect 23032 26382 23060 27270
rect 23020 26376 23072 26382
rect 23020 26318 23072 26324
rect 23124 25129 23152 28018
rect 23216 25498 23244 32932
rect 23492 32858 23520 33322
rect 23572 33108 23624 33114
rect 23572 33050 23624 33056
rect 23584 32978 23612 33050
rect 23572 32972 23624 32978
rect 23572 32914 23624 32920
rect 23296 32836 23348 32842
rect 23492 32830 23612 32858
rect 23296 32778 23348 32784
rect 23308 31414 23336 32778
rect 23480 31816 23532 31822
rect 23480 31758 23532 31764
rect 23296 31408 23348 31414
rect 23296 31350 23348 31356
rect 23296 31136 23348 31142
rect 23296 31078 23348 31084
rect 23308 30734 23336 31078
rect 23492 30870 23520 31758
rect 23480 30864 23532 30870
rect 23480 30806 23532 30812
rect 23492 30734 23520 30806
rect 23296 30728 23348 30734
rect 23296 30670 23348 30676
rect 23480 30728 23532 30734
rect 23480 30670 23532 30676
rect 23492 30394 23520 30670
rect 23480 30388 23532 30394
rect 23480 30330 23532 30336
rect 23584 30258 23612 32830
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23572 29232 23624 29238
rect 23572 29174 23624 29180
rect 23296 28960 23348 28966
rect 23296 28902 23348 28908
rect 23204 25492 23256 25498
rect 23204 25434 23256 25440
rect 23204 25220 23256 25226
rect 23204 25162 23256 25168
rect 23110 25120 23166 25129
rect 23110 25055 23166 25064
rect 23216 24834 23244 25162
rect 23124 24806 23244 24834
rect 22928 24608 22980 24614
rect 22926 24576 22928 24585
rect 22980 24576 22982 24585
rect 22926 24511 22982 24520
rect 22744 24404 22796 24410
rect 22744 24346 22796 24352
rect 22836 24404 22888 24410
rect 22836 24346 22888 24352
rect 22756 24138 22784 24346
rect 22744 24132 22796 24138
rect 22744 24074 22796 24080
rect 22664 22066 22784 22094
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22664 20806 22692 21966
rect 22652 20800 22704 20806
rect 22652 20742 22704 20748
rect 22664 20262 22692 20742
rect 22652 20256 22704 20262
rect 22652 20198 22704 20204
rect 22560 19712 22612 19718
rect 22560 19654 22612 19660
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22572 19378 22600 19654
rect 22664 19446 22692 19654
rect 22652 19440 22704 19446
rect 22652 19382 22704 19388
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22192 19168 22244 19174
rect 22192 19110 22244 19116
rect 22284 19168 22336 19174
rect 22284 19110 22336 19116
rect 22296 18986 22324 19110
rect 22204 18958 22324 18986
rect 22098 18456 22154 18465
rect 22098 18391 22100 18400
rect 22152 18391 22154 18400
rect 22100 18362 22152 18368
rect 22100 17672 22152 17678
rect 22100 17614 22152 17620
rect 22112 16726 22140 17614
rect 22100 16720 22152 16726
rect 22100 16662 22152 16668
rect 22112 16250 22140 16662
rect 22204 16538 22232 18958
rect 22468 18760 22520 18766
rect 22468 18702 22520 18708
rect 22480 17882 22508 18702
rect 22468 17876 22520 17882
rect 22468 17818 22520 17824
rect 22480 17678 22508 17818
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22284 17536 22336 17542
rect 22284 17478 22336 17484
rect 22468 17536 22520 17542
rect 22468 17478 22520 17484
rect 22296 16658 22324 17478
rect 22480 17202 22508 17478
rect 22468 17196 22520 17202
rect 22468 17138 22520 17144
rect 22466 17096 22522 17105
rect 22466 17031 22468 17040
rect 22520 17031 22522 17040
rect 22468 17002 22520 17008
rect 22376 16992 22428 16998
rect 22376 16934 22428 16940
rect 22388 16697 22416 16934
rect 22374 16688 22430 16697
rect 22284 16652 22336 16658
rect 22374 16623 22430 16632
rect 22468 16652 22520 16658
rect 22284 16594 22336 16600
rect 22468 16594 22520 16600
rect 22204 16510 22324 16538
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22204 16114 22232 16390
rect 22192 16108 22244 16114
rect 22192 16050 22244 16056
rect 22296 15994 22324 16510
rect 22204 15966 22324 15994
rect 22100 15428 22152 15434
rect 22100 15370 22152 15376
rect 22112 15162 22140 15370
rect 22100 15156 22152 15162
rect 22100 15098 22152 15104
rect 22100 12096 22152 12102
rect 22100 12038 22152 12044
rect 22112 11762 22140 12038
rect 22100 11756 22152 11762
rect 22100 11698 22152 11704
rect 22204 10010 22232 15966
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15026 22324 15846
rect 22480 15706 22508 16594
rect 22572 16522 22600 19314
rect 22652 18828 22704 18834
rect 22652 18770 22704 18776
rect 22664 17814 22692 18770
rect 22652 17808 22704 17814
rect 22652 17750 22704 17756
rect 22652 17604 22704 17610
rect 22652 17546 22704 17552
rect 22664 17513 22692 17546
rect 22650 17504 22706 17513
rect 22650 17439 22706 17448
rect 22652 17128 22704 17134
rect 22652 17070 22704 17076
rect 22664 16794 22692 17070
rect 22652 16788 22704 16794
rect 22652 16730 22704 16736
rect 22560 16516 22612 16522
rect 22560 16458 22612 16464
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 16114 22692 16390
rect 22652 16108 22704 16114
rect 22652 16050 22704 16056
rect 22468 15700 22520 15706
rect 22468 15642 22520 15648
rect 22480 15026 22508 15642
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 22468 15020 22520 15026
rect 22468 14962 22520 14968
rect 22652 12640 22704 12646
rect 22652 12582 22704 12588
rect 22664 12306 22692 12582
rect 22652 12300 22704 12306
rect 22652 12242 22704 12248
rect 22112 9982 22232 10010
rect 22112 8022 22140 9982
rect 22192 9920 22244 9926
rect 22192 9862 22244 9868
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 22204 7886 22232 9862
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22192 7880 22244 7886
rect 22192 7822 22244 7828
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22112 7154 22140 7754
rect 22204 7546 22232 7822
rect 22296 7818 22324 7958
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22284 7812 22336 7818
rect 22284 7754 22336 7760
rect 22192 7540 22244 7546
rect 22192 7482 22244 7488
rect 22112 7126 22232 7154
rect 22100 6996 22152 7002
rect 22100 6938 22152 6944
rect 22112 6390 22140 6938
rect 22204 6458 22232 7126
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 22296 6254 22324 7754
rect 22284 6248 22336 6254
rect 22284 6190 22336 6196
rect 22192 4548 22244 4554
rect 22192 4490 22244 4496
rect 22204 4282 22232 4490
rect 22192 4276 22244 4282
rect 22192 4218 22244 4224
rect 22560 4140 22612 4146
rect 22560 4082 22612 4088
rect 22468 4072 22520 4078
rect 22572 4049 22600 4082
rect 22468 4014 22520 4020
rect 22558 4040 22614 4049
rect 22480 3602 22508 4014
rect 22558 3975 22614 3984
rect 22664 3738 22692 7822
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22560 3052 22612 3058
rect 22560 2994 22612 3000
rect 21836 2746 22048 2774
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21272 2576 21324 2582
rect 21272 2518 21324 2524
rect 21180 2032 21232 2038
rect 21180 1974 21232 1980
rect 21284 800 21312 2518
rect 21836 2106 21864 2746
rect 21824 2100 21876 2106
rect 21824 2042 21876 2048
rect 22572 800 22600 2994
rect 22756 2854 22784 22066
rect 22848 14414 22876 24346
rect 23020 24336 23072 24342
rect 23020 24278 23072 24284
rect 23032 23798 23060 24278
rect 23020 23792 23072 23798
rect 23020 23734 23072 23740
rect 23020 23656 23072 23662
rect 23020 23598 23072 23604
rect 22928 23588 22980 23594
rect 22928 23530 22980 23536
rect 22940 23118 22968 23530
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 23032 22642 23060 23598
rect 23020 22636 23072 22642
rect 23020 22578 23072 22584
rect 22928 18148 22980 18154
rect 22928 18090 22980 18096
rect 22940 17746 22968 18090
rect 23020 17876 23072 17882
rect 23020 17818 23072 17824
rect 22928 17740 22980 17746
rect 22928 17682 22980 17688
rect 23032 17626 23060 17818
rect 22940 17598 23060 17626
rect 22940 17542 22968 17598
rect 22928 17536 22980 17542
rect 22928 17478 22980 17484
rect 23020 17536 23072 17542
rect 23020 17478 23072 17484
rect 22926 17368 22982 17377
rect 22926 17303 22982 17312
rect 22940 16658 22968 17303
rect 23032 16726 23060 17478
rect 23020 16720 23072 16726
rect 23020 16662 23072 16668
rect 22928 16652 22980 16658
rect 22928 16594 22980 16600
rect 22940 16153 22968 16594
rect 23020 16448 23072 16454
rect 23020 16390 23072 16396
rect 22926 16144 22982 16153
rect 23032 16114 23060 16390
rect 22926 16079 22982 16088
rect 23020 16108 23072 16114
rect 23020 16050 23072 16056
rect 22928 16040 22980 16046
rect 23124 15994 23152 24806
rect 23204 24608 23256 24614
rect 23204 24550 23256 24556
rect 23216 20369 23244 24550
rect 23308 23866 23336 28902
rect 23388 28552 23440 28558
rect 23388 28494 23440 28500
rect 23400 27033 23428 28494
rect 23584 28218 23612 29174
rect 23676 28490 23704 33476
rect 23848 33458 23900 33464
rect 23848 32496 23900 32502
rect 23848 32438 23900 32444
rect 23860 31278 23888 32438
rect 23848 31272 23900 31278
rect 23848 31214 23900 31220
rect 23756 29844 23808 29850
rect 23756 29786 23808 29792
rect 23768 29238 23796 29786
rect 23756 29232 23808 29238
rect 23756 29174 23808 29180
rect 23768 28762 23796 29174
rect 23756 28756 23808 28762
rect 23756 28698 23808 28704
rect 23664 28484 23716 28490
rect 23664 28426 23716 28432
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23664 28212 23716 28218
rect 23664 28154 23716 28160
rect 23676 27470 23704 28154
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23386 27024 23442 27033
rect 23386 26959 23442 26968
rect 23400 26246 23428 26959
rect 23676 26314 23704 27406
rect 23754 27296 23810 27305
rect 23754 27231 23810 27240
rect 23768 26926 23796 27231
rect 23952 26926 23980 34070
rect 24412 33862 24440 36042
rect 24504 35698 24532 39374
rect 24688 39370 24716 40870
rect 24676 39364 24728 39370
rect 24676 39306 24728 39312
rect 24688 38282 24716 39306
rect 24676 38276 24728 38282
rect 24676 38218 24728 38224
rect 24584 36848 24636 36854
rect 24584 36790 24636 36796
rect 24596 36582 24624 36790
rect 24584 36576 24636 36582
rect 24584 36518 24636 36524
rect 24584 36032 24636 36038
rect 24584 35974 24636 35980
rect 24492 35692 24544 35698
rect 24492 35634 24544 35640
rect 24504 35018 24532 35634
rect 24596 35630 24624 35974
rect 24676 35828 24728 35834
rect 24676 35770 24728 35776
rect 24584 35624 24636 35630
rect 24584 35566 24636 35572
rect 24584 35284 24636 35290
rect 24584 35226 24636 35232
rect 24596 35193 24624 35226
rect 24688 35222 24716 35770
rect 24676 35216 24728 35222
rect 24582 35184 24638 35193
rect 24676 35158 24728 35164
rect 24582 35119 24638 35128
rect 24492 35012 24544 35018
rect 24492 34954 24544 34960
rect 24596 34746 24624 35119
rect 24584 34740 24636 34746
rect 24584 34682 24636 34688
rect 24676 34672 24728 34678
rect 24676 34614 24728 34620
rect 24688 33930 24716 34614
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 24400 33856 24452 33862
rect 24400 33798 24452 33804
rect 24124 33652 24176 33658
rect 24124 33594 24176 33600
rect 24030 33552 24086 33561
rect 24030 33487 24032 33496
rect 24084 33487 24086 33496
rect 24032 33458 24084 33464
rect 24032 33312 24084 33318
rect 24032 33254 24084 33260
rect 24044 32434 24072 33254
rect 24032 32428 24084 32434
rect 24032 32370 24084 32376
rect 24032 31340 24084 31346
rect 24032 31282 24084 31288
rect 24044 28490 24072 31282
rect 24032 28484 24084 28490
rect 24032 28426 24084 28432
rect 24044 28150 24072 28426
rect 24032 28144 24084 28150
rect 24032 28086 24084 28092
rect 23756 26920 23808 26926
rect 23756 26862 23808 26868
rect 23940 26920 23992 26926
rect 23940 26862 23992 26868
rect 24032 26512 24084 26518
rect 24032 26454 24084 26460
rect 23664 26308 23716 26314
rect 23664 26250 23716 26256
rect 24044 26246 24072 26454
rect 23388 26240 23440 26246
rect 23388 26182 23440 26188
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 23400 24614 23428 26182
rect 23480 25900 23532 25906
rect 23480 25842 23532 25848
rect 23492 25378 23520 25842
rect 23572 25832 23624 25838
rect 23572 25774 23624 25780
rect 23584 25498 23612 25774
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23572 25492 23624 25498
rect 23572 25434 23624 25440
rect 23492 25350 23704 25378
rect 23676 25106 23704 25350
rect 23492 25078 23704 25106
rect 23492 24954 23520 25078
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23388 24608 23440 24614
rect 23388 24550 23440 24556
rect 23664 24608 23716 24614
rect 23664 24550 23716 24556
rect 23296 23860 23348 23866
rect 23296 23802 23348 23808
rect 23308 23118 23336 23802
rect 23676 23780 23704 24550
rect 23584 23752 23704 23780
rect 23296 23112 23348 23118
rect 23296 23054 23348 23060
rect 23584 22982 23612 23752
rect 23768 23662 23796 24754
rect 23952 24274 23980 25638
rect 24032 24880 24084 24886
rect 24032 24822 24084 24828
rect 23940 24268 23992 24274
rect 23940 24210 23992 24216
rect 23846 24168 23902 24177
rect 23846 24103 23902 24112
rect 23860 23730 23888 24103
rect 23848 23724 23900 23730
rect 23848 23666 23900 23672
rect 23756 23656 23808 23662
rect 23756 23598 23808 23604
rect 23664 23520 23716 23526
rect 23664 23462 23716 23468
rect 23572 22976 23624 22982
rect 23572 22918 23624 22924
rect 23570 22536 23626 22545
rect 23570 22471 23626 22480
rect 23480 21344 23532 21350
rect 23480 21286 23532 21292
rect 23492 20942 23520 21286
rect 23480 20936 23532 20942
rect 23480 20878 23532 20884
rect 23480 20596 23532 20602
rect 23480 20538 23532 20544
rect 23294 20496 23350 20505
rect 23492 20466 23520 20538
rect 23294 20431 23296 20440
rect 23348 20431 23350 20440
rect 23480 20460 23532 20466
rect 23296 20402 23348 20408
rect 23480 20402 23532 20408
rect 23202 20360 23258 20369
rect 23202 20295 23258 20304
rect 23204 20256 23256 20262
rect 23204 20198 23256 20204
rect 23216 19446 23244 20198
rect 23204 19440 23256 19446
rect 23204 19382 23256 19388
rect 23204 18284 23256 18290
rect 23204 18226 23256 18232
rect 23480 18284 23532 18290
rect 23480 18226 23532 18232
rect 23216 17202 23244 18226
rect 23296 18080 23348 18086
rect 23296 18022 23348 18028
rect 23308 17678 23336 18022
rect 23492 17814 23520 18226
rect 23480 17808 23532 17814
rect 23480 17750 23532 17756
rect 23388 17740 23440 17746
rect 23388 17682 23440 17688
rect 23296 17672 23348 17678
rect 23400 17649 23428 17682
rect 23296 17614 23348 17620
rect 23386 17640 23442 17649
rect 23308 17270 23336 17614
rect 23386 17575 23442 17584
rect 23386 17504 23442 17513
rect 23386 17439 23442 17448
rect 23400 17270 23428 17439
rect 23296 17264 23348 17270
rect 23296 17206 23348 17212
rect 23388 17264 23440 17270
rect 23388 17206 23440 17212
rect 23204 17196 23256 17202
rect 23204 17138 23256 17144
rect 23388 17128 23440 17134
rect 23388 17070 23440 17076
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23308 16708 23336 17002
rect 23400 16833 23428 17070
rect 23386 16824 23442 16833
rect 23386 16759 23442 16768
rect 23308 16680 23428 16708
rect 23296 16516 23348 16522
rect 23296 16458 23348 16464
rect 22928 15982 22980 15988
rect 22940 15706 22968 15982
rect 23032 15966 23152 15994
rect 22928 15700 22980 15706
rect 22928 15642 22980 15648
rect 22836 14408 22888 14414
rect 22836 14350 22888 14356
rect 22836 12096 22888 12102
rect 22836 12038 22888 12044
rect 22848 11694 22876 12038
rect 22836 11688 22888 11694
rect 22836 11630 22888 11636
rect 22848 11354 22876 11630
rect 22836 11348 22888 11354
rect 22836 11290 22888 11296
rect 22744 2848 22796 2854
rect 22744 2790 22796 2796
rect 23032 2310 23060 15966
rect 23308 15502 23336 16458
rect 23400 16402 23428 16680
rect 23492 16658 23520 17750
rect 23480 16652 23532 16658
rect 23480 16594 23532 16600
rect 23478 16552 23534 16561
rect 23478 16487 23480 16496
rect 23532 16487 23534 16496
rect 23480 16458 23532 16464
rect 23400 16374 23520 16402
rect 23112 15496 23164 15502
rect 23112 15438 23164 15444
rect 23296 15496 23348 15502
rect 23296 15438 23348 15444
rect 23124 15094 23152 15438
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23492 14822 23520 16374
rect 23388 14816 23440 14822
rect 23388 14758 23440 14764
rect 23480 14816 23532 14822
rect 23480 14758 23532 14764
rect 23400 14634 23428 14758
rect 23400 14618 23520 14634
rect 23400 14612 23532 14618
rect 23400 14606 23480 14612
rect 23480 14554 23532 14560
rect 23296 13728 23348 13734
rect 23296 13670 23348 13676
rect 23308 13326 23336 13670
rect 23480 13388 23532 13394
rect 23480 13330 23532 13336
rect 23296 13320 23348 13326
rect 23296 13262 23348 13268
rect 23388 13184 23440 13190
rect 23388 13126 23440 13132
rect 23204 12844 23256 12850
rect 23204 12786 23256 12792
rect 23296 12844 23348 12850
rect 23296 12786 23348 12792
rect 23216 11762 23244 12786
rect 23204 11756 23256 11762
rect 23204 11698 23256 11704
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 23124 10062 23152 10542
rect 23112 10056 23164 10062
rect 23112 9998 23164 10004
rect 23308 9926 23336 12786
rect 23400 12102 23428 13126
rect 23492 12986 23520 13330
rect 23480 12980 23532 12986
rect 23480 12922 23532 12928
rect 23480 12708 23532 12714
rect 23480 12650 23532 12656
rect 23388 12096 23440 12102
rect 23388 12038 23440 12044
rect 23492 11898 23520 12650
rect 23480 11892 23532 11898
rect 23480 11834 23532 11840
rect 23480 10532 23532 10538
rect 23480 10474 23532 10480
rect 23492 10266 23520 10474
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23480 10056 23532 10062
rect 23480 9998 23532 10004
rect 23492 9926 23520 9998
rect 23296 9920 23348 9926
rect 23296 9862 23348 9868
rect 23480 9920 23532 9926
rect 23480 9862 23532 9868
rect 23584 7970 23612 22471
rect 23676 21554 23704 23462
rect 23768 22234 23796 23598
rect 23860 22710 23888 23666
rect 23940 23316 23992 23322
rect 23940 23258 23992 23264
rect 23848 22704 23900 22710
rect 23848 22646 23900 22652
rect 23952 22506 23980 23258
rect 24044 23186 24072 24822
rect 24136 24750 24164 33594
rect 24308 33448 24360 33454
rect 24308 33390 24360 33396
rect 24320 33114 24348 33390
rect 24308 33108 24360 33114
rect 24308 33050 24360 33056
rect 24308 32972 24360 32978
rect 24308 32914 24360 32920
rect 24320 31482 24348 32914
rect 24308 31476 24360 31482
rect 24308 31418 24360 31424
rect 24320 30870 24348 31418
rect 24412 31346 24440 33798
rect 24688 32978 24716 33866
rect 24676 32972 24728 32978
rect 24676 32914 24728 32920
rect 24780 31754 24808 46582
rect 24860 40452 24912 40458
rect 24860 40394 24912 40400
rect 24872 39846 24900 40394
rect 25320 40112 25372 40118
rect 25320 40054 25372 40060
rect 25044 40044 25096 40050
rect 25044 39986 25096 39992
rect 24952 39908 25004 39914
rect 24952 39850 25004 39856
rect 24860 39840 24912 39846
rect 24860 39782 24912 39788
rect 24872 38570 24900 39782
rect 24964 39030 24992 39850
rect 25056 39098 25084 39986
rect 25136 39296 25188 39302
rect 25136 39238 25188 39244
rect 25044 39092 25096 39098
rect 25044 39034 25096 39040
rect 25148 39030 25176 39238
rect 24952 39024 25004 39030
rect 24952 38966 25004 38972
rect 25136 39024 25188 39030
rect 25136 38966 25188 38972
rect 24964 38758 24992 38966
rect 25228 38888 25280 38894
rect 25228 38830 25280 38836
rect 24952 38752 25004 38758
rect 24952 38694 25004 38700
rect 25136 38752 25188 38758
rect 25136 38694 25188 38700
rect 24872 38542 25084 38570
rect 24952 38344 25004 38350
rect 24952 38286 25004 38292
rect 24964 38010 24992 38286
rect 25056 38196 25084 38542
rect 25148 38350 25176 38694
rect 25136 38344 25188 38350
rect 25136 38286 25188 38292
rect 25056 38168 25176 38196
rect 24860 38004 24912 38010
rect 24860 37946 24912 37952
rect 24952 38004 25004 38010
rect 24952 37946 25004 37952
rect 24872 34066 24900 37946
rect 25148 37874 25176 38168
rect 25136 37868 25188 37874
rect 25136 37810 25188 37816
rect 24952 37800 25004 37806
rect 24952 37742 25004 37748
rect 24964 37330 24992 37742
rect 24952 37324 25004 37330
rect 24952 37266 25004 37272
rect 25148 35018 25176 37810
rect 25136 35012 25188 35018
rect 25136 34954 25188 34960
rect 25136 34400 25188 34406
rect 25136 34342 25188 34348
rect 24860 34060 24912 34066
rect 24860 34002 24912 34008
rect 24872 33946 24900 34002
rect 25148 33998 25176 34342
rect 25136 33992 25188 33998
rect 24872 33918 24992 33946
rect 25136 33934 25188 33940
rect 24964 32994 24992 33918
rect 25136 33584 25188 33590
rect 25136 33526 25188 33532
rect 25044 33380 25096 33386
rect 25044 33322 25096 33328
rect 24688 31726 24808 31754
rect 24872 32966 24992 32994
rect 24400 31340 24452 31346
rect 24400 31282 24452 31288
rect 24308 30864 24360 30870
rect 24308 30806 24360 30812
rect 24308 30592 24360 30598
rect 24308 30534 24360 30540
rect 24320 30054 24348 30534
rect 24308 30048 24360 30054
rect 24308 29990 24360 29996
rect 24320 29510 24348 29990
rect 24308 29504 24360 29510
rect 24308 29446 24360 29452
rect 24584 25900 24636 25906
rect 24584 25842 24636 25848
rect 24492 25424 24544 25430
rect 24492 25366 24544 25372
rect 24504 25129 24532 25366
rect 24596 25294 24624 25842
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24490 25120 24546 25129
rect 24490 25055 24546 25064
rect 24688 24993 24716 31726
rect 24768 31408 24820 31414
rect 24768 31350 24820 31356
rect 24780 30938 24808 31350
rect 24768 30932 24820 30938
rect 24768 30874 24820 30880
rect 24780 28762 24808 30874
rect 24872 30802 24900 32966
rect 24952 32564 25004 32570
rect 24952 32506 25004 32512
rect 24964 32366 24992 32506
rect 24952 32360 25004 32366
rect 24952 32302 25004 32308
rect 25056 32178 25084 33322
rect 24964 32150 25084 32178
rect 24860 30796 24912 30802
rect 24860 30738 24912 30744
rect 24964 30394 24992 32150
rect 25148 31754 25176 33526
rect 25240 32042 25268 38830
rect 25332 38486 25360 40054
rect 25320 38480 25372 38486
rect 25320 38422 25372 38428
rect 25332 37738 25360 38422
rect 25320 37732 25372 37738
rect 25320 37674 25372 37680
rect 25320 34604 25372 34610
rect 25320 34546 25372 34552
rect 25332 32570 25360 34546
rect 25424 34082 25452 49030
rect 26700 48544 26752 48550
rect 26700 48486 26752 48492
rect 26712 48210 26740 48486
rect 27080 48210 27108 51200
rect 27712 49156 27764 49162
rect 27712 49098 27764 49104
rect 27252 48680 27304 48686
rect 27252 48622 27304 48628
rect 26700 48204 26752 48210
rect 26700 48146 26752 48152
rect 27068 48204 27120 48210
rect 27068 48146 27120 48152
rect 26332 48068 26384 48074
rect 26332 48010 26384 48016
rect 26344 47802 26372 48010
rect 27264 47802 27292 48622
rect 26332 47796 26384 47802
rect 26332 47738 26384 47744
rect 27252 47796 27304 47802
rect 27252 47738 27304 47744
rect 26516 47728 26568 47734
rect 26516 47670 26568 47676
rect 26424 47592 26476 47598
rect 26424 47534 26476 47540
rect 26436 45830 26464 47534
rect 26424 45824 26476 45830
rect 26424 45766 26476 45772
rect 25872 42152 25924 42158
rect 25872 42094 25924 42100
rect 25884 40050 25912 42094
rect 25872 40044 25924 40050
rect 25872 39986 25924 39992
rect 25780 39976 25832 39982
rect 25780 39918 25832 39924
rect 25688 39364 25740 39370
rect 25688 39306 25740 39312
rect 25700 39098 25728 39306
rect 25792 39302 25820 39918
rect 26148 39840 26200 39846
rect 26148 39782 26200 39788
rect 26056 39500 26108 39506
rect 26056 39442 26108 39448
rect 25780 39296 25832 39302
rect 25780 39238 25832 39244
rect 25688 39092 25740 39098
rect 25688 39034 25740 39040
rect 25792 38962 25820 39238
rect 25780 38956 25832 38962
rect 25780 38898 25832 38904
rect 26068 38758 26096 39442
rect 26160 38962 26188 39782
rect 26148 38956 26200 38962
rect 26148 38898 26200 38904
rect 26056 38752 26108 38758
rect 26056 38694 26108 38700
rect 25688 38208 25740 38214
rect 25688 38150 25740 38156
rect 25700 35154 25728 38150
rect 25780 37868 25832 37874
rect 25780 37810 25832 37816
rect 25792 37194 25820 37810
rect 25780 37188 25832 37194
rect 25780 37130 25832 37136
rect 25792 36922 25820 37130
rect 25872 37120 25924 37126
rect 25872 37062 25924 37068
rect 25780 36916 25832 36922
rect 25780 36858 25832 36864
rect 25884 36786 25912 37062
rect 25872 36780 25924 36786
rect 25872 36722 25924 36728
rect 25780 35828 25832 35834
rect 25780 35770 25832 35776
rect 25504 35148 25556 35154
rect 25504 35090 25556 35096
rect 25688 35148 25740 35154
rect 25688 35090 25740 35096
rect 25516 34202 25544 35090
rect 25596 34944 25648 34950
rect 25596 34886 25648 34892
rect 25504 34196 25556 34202
rect 25504 34138 25556 34144
rect 25424 34054 25544 34082
rect 25410 33552 25466 33561
rect 25410 33487 25412 33496
rect 25464 33487 25466 33496
rect 25412 33458 25464 33464
rect 25320 32564 25372 32570
rect 25320 32506 25372 32512
rect 25332 32230 25360 32506
rect 25320 32224 25372 32230
rect 25320 32166 25372 32172
rect 25240 32014 25360 32042
rect 25228 31816 25280 31822
rect 25228 31758 25280 31764
rect 25136 31748 25188 31754
rect 25136 31690 25188 31696
rect 25044 31272 25096 31278
rect 25044 31214 25096 31220
rect 24952 30388 25004 30394
rect 24952 30330 25004 30336
rect 25056 30258 25084 31214
rect 25148 30666 25176 31690
rect 25136 30660 25188 30666
rect 25136 30602 25188 30608
rect 25044 30252 25096 30258
rect 25096 30212 25176 30240
rect 25044 30194 25096 30200
rect 25044 30048 25096 30054
rect 25044 29990 25096 29996
rect 25056 29034 25084 29990
rect 25044 29028 25096 29034
rect 25044 28970 25096 28976
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 25148 28558 25176 30212
rect 25136 28552 25188 28558
rect 25136 28494 25188 28500
rect 24952 28416 25004 28422
rect 24952 28358 25004 28364
rect 24860 28008 24912 28014
rect 24860 27950 24912 27956
rect 24872 26602 24900 27950
rect 24964 27674 24992 28358
rect 25148 28150 25176 28494
rect 25136 28144 25188 28150
rect 25136 28086 25188 28092
rect 24952 27668 25004 27674
rect 24952 27610 25004 27616
rect 24952 27464 25004 27470
rect 24952 27406 25004 27412
rect 24964 27130 24992 27406
rect 24952 27124 25004 27130
rect 24952 27066 25004 27072
rect 25044 27124 25096 27130
rect 25044 27066 25096 27072
rect 25056 26874 25084 27066
rect 24964 26846 25084 26874
rect 24964 26790 24992 26846
rect 24952 26784 25004 26790
rect 24952 26726 25004 26732
rect 24872 26574 24992 26602
rect 24964 26314 24992 26574
rect 25240 26518 25268 31758
rect 25332 28994 25360 32014
rect 25516 30870 25544 34054
rect 25504 30864 25556 30870
rect 25504 30806 25556 30812
rect 25608 30682 25636 34886
rect 25792 32994 25820 35770
rect 25884 34406 25912 36722
rect 25964 36576 26016 36582
rect 25964 36518 26016 36524
rect 25976 36106 26004 36518
rect 25964 36100 26016 36106
rect 25964 36042 26016 36048
rect 25872 34400 25924 34406
rect 25872 34342 25924 34348
rect 26068 34354 26096 38694
rect 26240 37664 26292 37670
rect 26240 37606 26292 37612
rect 26252 37398 26280 37606
rect 26240 37392 26292 37398
rect 26240 37334 26292 37340
rect 26148 37324 26200 37330
rect 26148 37266 26200 37272
rect 26160 36718 26188 37266
rect 26148 36712 26200 36718
rect 26148 36654 26200 36660
rect 26160 35578 26188 36654
rect 26332 36576 26384 36582
rect 26332 36518 26384 36524
rect 26344 36174 26372 36518
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26240 35624 26292 35630
rect 26238 35592 26240 35601
rect 26292 35592 26294 35601
rect 26160 35550 26238 35578
rect 26160 34542 26188 35550
rect 26238 35527 26294 35536
rect 26240 35080 26292 35086
rect 26240 35022 26292 35028
rect 26148 34536 26200 34542
rect 26148 34478 26200 34484
rect 26068 34326 26188 34354
rect 25964 34196 26016 34202
rect 25964 34138 26016 34144
rect 25976 33318 26004 34138
rect 25872 33312 25924 33318
rect 25872 33254 25924 33260
rect 25964 33312 26016 33318
rect 25964 33254 26016 33260
rect 25700 32966 25820 32994
rect 25700 32434 25728 32966
rect 25884 32910 25912 33254
rect 25780 32904 25832 32910
rect 25780 32846 25832 32852
rect 25872 32904 25924 32910
rect 25872 32846 25924 32852
rect 25792 32502 25820 32846
rect 25976 32774 26004 33254
rect 25964 32768 26016 32774
rect 25964 32710 26016 32716
rect 25780 32496 25832 32502
rect 25780 32438 25832 32444
rect 25688 32428 25740 32434
rect 25688 32370 25740 32376
rect 25700 32026 25728 32370
rect 25688 32020 25740 32026
rect 25688 31962 25740 31968
rect 25792 31686 25820 32438
rect 26160 32416 26188 34326
rect 26252 34202 26280 35022
rect 26240 34196 26292 34202
rect 26240 34138 26292 34144
rect 26332 34060 26384 34066
rect 26332 34002 26384 34008
rect 26344 32570 26372 34002
rect 26332 32564 26384 32570
rect 26332 32506 26384 32512
rect 26240 32428 26292 32434
rect 26160 32388 26240 32416
rect 26240 32370 26292 32376
rect 26148 32224 26200 32230
rect 26148 32166 26200 32172
rect 25780 31680 25832 31686
rect 25780 31622 25832 31628
rect 26160 31278 26188 32166
rect 26252 31822 26280 32370
rect 26332 31884 26384 31890
rect 26332 31826 26384 31832
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 26240 31408 26292 31414
rect 26240 31350 26292 31356
rect 26148 31272 26200 31278
rect 26148 31214 26200 31220
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25976 30870 26004 31078
rect 25872 30864 25924 30870
rect 25778 30832 25834 30841
rect 25872 30806 25924 30812
rect 25964 30864 26016 30870
rect 25964 30806 26016 30812
rect 25778 30767 25834 30776
rect 25792 30734 25820 30767
rect 25516 30654 25636 30682
rect 25780 30728 25832 30734
rect 25780 30670 25832 30676
rect 25412 30252 25464 30258
rect 25412 30194 25464 30200
rect 25424 29850 25452 30194
rect 25412 29844 25464 29850
rect 25412 29786 25464 29792
rect 25332 28966 25452 28994
rect 25320 27872 25372 27878
rect 25320 27814 25372 27820
rect 25332 27062 25360 27814
rect 25320 27056 25372 27062
rect 25320 26998 25372 27004
rect 25228 26512 25280 26518
rect 25056 26460 25228 26466
rect 25056 26454 25280 26460
rect 25056 26438 25268 26454
rect 24768 26308 24820 26314
rect 24768 26250 24820 26256
rect 24952 26308 25004 26314
rect 24952 26250 25004 26256
rect 24674 24984 24730 24993
rect 24674 24919 24730 24928
rect 24124 24744 24176 24750
rect 24124 24686 24176 24692
rect 24780 24614 24808 26250
rect 24860 25764 24912 25770
rect 24860 25706 24912 25712
rect 24872 25430 24900 25706
rect 24860 25424 24912 25430
rect 24860 25366 24912 25372
rect 24768 24608 24820 24614
rect 24214 24576 24270 24585
rect 24768 24550 24820 24556
rect 24214 24511 24270 24520
rect 24032 23180 24084 23186
rect 24032 23122 24084 23128
rect 24228 23066 24256 24511
rect 24308 24404 24360 24410
rect 24308 24346 24360 24352
rect 24320 23322 24348 24346
rect 24492 24268 24544 24274
rect 24492 24210 24544 24216
rect 24400 24200 24452 24206
rect 24400 24142 24452 24148
rect 24412 23730 24440 24142
rect 24400 23724 24452 23730
rect 24400 23666 24452 23672
rect 24308 23316 24360 23322
rect 24308 23258 24360 23264
rect 24228 23038 24348 23066
rect 24412 23050 24440 23666
rect 24504 23186 24532 24210
rect 24676 24200 24728 24206
rect 24674 24168 24676 24177
rect 24728 24168 24730 24177
rect 24674 24103 24730 24112
rect 24582 24032 24638 24041
rect 24582 23967 24638 23976
rect 24492 23180 24544 23186
rect 24492 23122 24544 23128
rect 24216 22976 24268 22982
rect 24216 22918 24268 22924
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 23756 22228 23808 22234
rect 23756 22170 23808 22176
rect 23952 22094 23980 22442
rect 23860 22066 23980 22094
rect 23860 22030 23888 22066
rect 23848 22024 23900 22030
rect 23848 21966 23900 21972
rect 23756 21956 23808 21962
rect 23756 21898 23808 21904
rect 23664 21548 23716 21554
rect 23664 21490 23716 21496
rect 23676 19718 23704 21490
rect 23664 19712 23716 19718
rect 23664 19654 23716 19660
rect 23664 18624 23716 18630
rect 23664 18566 23716 18572
rect 23676 17202 23704 18566
rect 23664 17196 23716 17202
rect 23664 17138 23716 17144
rect 23662 17096 23718 17105
rect 23662 17031 23664 17040
rect 23716 17031 23718 17040
rect 23664 17002 23716 17008
rect 23662 16144 23718 16153
rect 23662 16079 23664 16088
rect 23716 16079 23718 16088
rect 23664 16050 23716 16056
rect 23664 14816 23716 14822
rect 23664 14758 23716 14764
rect 23676 13870 23704 14758
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23676 12238 23704 12582
rect 23664 12232 23716 12238
rect 23664 12174 23716 12180
rect 23492 7942 23612 7970
rect 23664 8016 23716 8022
rect 23664 7958 23716 7964
rect 23388 6792 23440 6798
rect 23388 6734 23440 6740
rect 23400 6322 23428 6734
rect 23388 6316 23440 6322
rect 23388 6258 23440 6264
rect 23492 5914 23520 7942
rect 23676 7868 23704 7958
rect 23584 7840 23704 7868
rect 23584 6798 23612 7840
rect 23768 7562 23796 21898
rect 24124 21548 24176 21554
rect 24124 21490 24176 21496
rect 24032 21480 24084 21486
rect 24032 21422 24084 21428
rect 24044 20874 24072 21422
rect 24032 20868 24084 20874
rect 24032 20810 24084 20816
rect 23940 20392 23992 20398
rect 23940 20334 23992 20340
rect 23952 19446 23980 20334
rect 24044 20262 24072 20810
rect 24032 20256 24084 20262
rect 24032 20198 24084 20204
rect 23940 19440 23992 19446
rect 23940 19382 23992 19388
rect 23940 19304 23992 19310
rect 23940 19246 23992 19252
rect 24032 19304 24084 19310
rect 24032 19246 24084 19252
rect 23848 18080 23900 18086
rect 23848 18022 23900 18028
rect 23860 16794 23888 18022
rect 23848 16788 23900 16794
rect 23848 16730 23900 16736
rect 23846 16688 23902 16697
rect 23846 16623 23902 16632
rect 23860 14822 23888 16623
rect 23848 14816 23900 14822
rect 23848 14758 23900 14764
rect 23860 14006 23888 14758
rect 23848 14000 23900 14006
rect 23848 13942 23900 13948
rect 23848 13524 23900 13530
rect 23848 13466 23900 13472
rect 23860 12782 23888 13466
rect 23848 12776 23900 12782
rect 23848 12718 23900 12724
rect 23848 9920 23900 9926
rect 23848 9862 23900 9868
rect 23860 9586 23888 9862
rect 23848 9580 23900 9586
rect 23848 9522 23900 9528
rect 23848 8084 23900 8090
rect 23848 8026 23900 8032
rect 23860 7886 23888 8026
rect 23952 7970 23980 19246
rect 24044 18222 24072 19246
rect 24032 18216 24084 18222
rect 24032 18158 24084 18164
rect 24032 18080 24084 18086
rect 24032 18022 24084 18028
rect 24044 17202 24072 18022
rect 24136 17882 24164 21490
rect 24124 17876 24176 17882
rect 24124 17818 24176 17824
rect 24228 17218 24256 22918
rect 24320 20618 24348 23038
rect 24400 23044 24452 23050
rect 24400 22986 24452 22992
rect 24398 22944 24454 22953
rect 24398 22879 24454 22888
rect 24412 22234 24440 22879
rect 24400 22228 24452 22234
rect 24400 22170 24452 22176
rect 24504 22166 24532 23122
rect 24596 23118 24624 23967
rect 24676 23588 24728 23594
rect 24676 23530 24728 23536
rect 24584 23112 24636 23118
rect 24584 23054 24636 23060
rect 24596 22642 24624 23054
rect 24688 22710 24716 23530
rect 24676 22704 24728 22710
rect 24676 22646 24728 22652
rect 24584 22636 24636 22642
rect 24584 22578 24636 22584
rect 24492 22160 24544 22166
rect 24492 22102 24544 22108
rect 24400 21956 24452 21962
rect 24400 21898 24452 21904
rect 24412 20777 24440 21898
rect 24584 21888 24636 21894
rect 24582 21856 24584 21865
rect 24636 21856 24638 21865
rect 24582 21791 24638 21800
rect 24582 21720 24638 21729
rect 24582 21655 24638 21664
rect 24596 21418 24624 21655
rect 24584 21412 24636 21418
rect 24584 21354 24636 21360
rect 24492 21344 24544 21350
rect 24492 21286 24544 21292
rect 24504 20942 24532 21286
rect 24492 20936 24544 20942
rect 24492 20878 24544 20884
rect 24398 20768 24454 20777
rect 24398 20703 24454 20712
rect 24320 20590 24440 20618
rect 24308 20256 24360 20262
rect 24308 20198 24360 20204
rect 24032 17196 24084 17202
rect 24032 17138 24084 17144
rect 24136 17190 24256 17218
rect 24032 16176 24084 16182
rect 24032 16118 24084 16124
rect 24044 15026 24072 16118
rect 24136 15978 24164 17190
rect 24216 17060 24268 17066
rect 24216 17002 24268 17008
rect 24124 15972 24176 15978
rect 24124 15914 24176 15920
rect 24136 15434 24164 15914
rect 24124 15428 24176 15434
rect 24124 15370 24176 15376
rect 24032 15020 24084 15026
rect 24032 14962 24084 14968
rect 24124 13864 24176 13870
rect 24124 13806 24176 13812
rect 24032 13796 24084 13802
rect 24032 13738 24084 13744
rect 24044 12850 24072 13738
rect 24136 13190 24164 13806
rect 24124 13184 24176 13190
rect 24124 13126 24176 13132
rect 24032 12844 24084 12850
rect 24032 12786 24084 12792
rect 24136 12782 24164 13126
rect 24124 12776 24176 12782
rect 24124 12718 24176 12724
rect 24032 12232 24084 12238
rect 24032 12174 24084 12180
rect 24044 10674 24072 12174
rect 24136 11150 24164 12718
rect 24124 11144 24176 11150
rect 24124 11086 24176 11092
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 10266 24072 10610
rect 24032 10260 24084 10266
rect 24032 10202 24084 10208
rect 23952 7942 24164 7970
rect 23848 7880 23900 7886
rect 23900 7840 24072 7868
rect 23848 7822 23900 7828
rect 23768 7534 23980 7562
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23768 6866 23796 7346
rect 23756 6860 23808 6866
rect 23756 6802 23808 6808
rect 23572 6792 23624 6798
rect 23572 6734 23624 6740
rect 23664 6792 23716 6798
rect 23664 6734 23716 6740
rect 23584 6662 23612 6734
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23676 6458 23704 6734
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23296 3732 23348 3738
rect 23296 3674 23348 3680
rect 23308 3534 23336 3674
rect 23204 3528 23256 3534
rect 23204 3470 23256 3476
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23020 2304 23072 2310
rect 23020 2246 23072 2252
rect 23216 800 23244 3470
rect 23308 3126 23336 3470
rect 23296 3120 23348 3126
rect 23296 3062 23348 3068
rect 23400 3058 23428 3878
rect 23572 3392 23624 3398
rect 23572 3334 23624 3340
rect 23584 3126 23612 3334
rect 23572 3120 23624 3126
rect 23572 3062 23624 3068
rect 23388 3052 23440 3058
rect 23388 2994 23440 3000
rect 23848 2984 23900 2990
rect 23848 2926 23900 2932
rect 23860 800 23888 2926
rect 23952 2514 23980 7534
rect 24044 6798 24072 7840
rect 24032 6792 24084 6798
rect 24032 6734 24084 6740
rect 24136 2990 24164 7942
rect 24124 2984 24176 2990
rect 24124 2926 24176 2932
rect 24228 2774 24256 17002
rect 24320 13530 24348 20198
rect 24412 18630 24440 20590
rect 24688 19258 24716 22646
rect 24780 21486 24808 24550
rect 24860 22636 24912 22642
rect 24860 22578 24912 22584
rect 24768 21480 24820 21486
rect 24768 21422 24820 21428
rect 24768 19712 24820 19718
rect 24768 19654 24820 19660
rect 24504 19230 24716 19258
rect 24400 18624 24452 18630
rect 24400 18566 24452 18572
rect 24504 16674 24532 19230
rect 24676 19168 24728 19174
rect 24676 19110 24728 19116
rect 24688 18766 24716 19110
rect 24676 18760 24728 18766
rect 24676 18702 24728 18708
rect 24584 18624 24636 18630
rect 24584 18566 24636 18572
rect 24596 17898 24624 18566
rect 24688 18426 24716 18702
rect 24676 18420 24728 18426
rect 24676 18362 24728 18368
rect 24688 18154 24716 18362
rect 24676 18148 24728 18154
rect 24676 18090 24728 18096
rect 24596 17870 24716 17898
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24596 17134 24624 17546
rect 24584 17128 24636 17134
rect 24584 17070 24636 17076
rect 24504 16646 24624 16674
rect 24492 16516 24544 16522
rect 24492 16458 24544 16464
rect 24400 16448 24452 16454
rect 24400 16390 24452 16396
rect 24412 16250 24440 16390
rect 24400 16244 24452 16250
rect 24400 16186 24452 16192
rect 24504 15502 24532 16458
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24596 15314 24624 16646
rect 24688 16182 24716 17870
rect 24676 16176 24728 16182
rect 24676 16118 24728 16124
rect 24504 15286 24624 15314
rect 24400 15020 24452 15026
rect 24400 14962 24452 14968
rect 24308 13524 24360 13530
rect 24308 13466 24360 13472
rect 24412 12850 24440 14962
rect 24504 14618 24532 15286
rect 24688 15144 24716 16118
rect 24780 15706 24808 19654
rect 24872 17338 24900 22578
rect 24964 18766 24992 26250
rect 24952 18760 25004 18766
rect 24952 18702 25004 18708
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 24964 17814 24992 18226
rect 24952 17808 25004 17814
rect 24952 17750 25004 17756
rect 24952 17536 25004 17542
rect 24952 17478 25004 17484
rect 24860 17332 24912 17338
rect 24860 17274 24912 17280
rect 24860 16720 24912 16726
rect 24860 16662 24912 16668
rect 24872 16046 24900 16662
rect 24964 16182 24992 17478
rect 24952 16176 25004 16182
rect 24952 16118 25004 16124
rect 24860 16040 24912 16046
rect 24860 15982 24912 15988
rect 24768 15700 24820 15706
rect 24768 15642 24820 15648
rect 24596 15116 24716 15144
rect 24596 15026 24624 15116
rect 24780 15042 24808 15642
rect 24584 15020 24636 15026
rect 24584 14962 24636 14968
rect 24688 15014 24808 15042
rect 24872 15026 24900 15982
rect 24964 15502 24992 16118
rect 25056 16114 25084 26438
rect 25228 26036 25280 26042
rect 25228 25978 25280 25984
rect 25136 25832 25188 25838
rect 25136 25774 25188 25780
rect 25148 25498 25176 25774
rect 25240 25770 25268 25978
rect 25228 25764 25280 25770
rect 25228 25706 25280 25712
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25136 22636 25188 22642
rect 25136 22578 25188 22584
rect 25148 22234 25176 22578
rect 25320 22568 25372 22574
rect 25320 22510 25372 22516
rect 25228 22432 25280 22438
rect 25228 22374 25280 22380
rect 25136 22228 25188 22234
rect 25136 22170 25188 22176
rect 25240 22094 25268 22374
rect 25148 22066 25268 22094
rect 25148 21146 25176 22066
rect 25228 22024 25280 22030
rect 25228 21966 25280 21972
rect 25136 21140 25188 21146
rect 25136 21082 25188 21088
rect 25136 18692 25188 18698
rect 25136 18634 25188 18640
rect 25148 17678 25176 18634
rect 25136 17672 25188 17678
rect 25136 17614 25188 17620
rect 25136 16788 25188 16794
rect 25136 16730 25188 16736
rect 25044 16108 25096 16114
rect 25044 16050 25096 16056
rect 24952 15496 25004 15502
rect 24952 15438 25004 15444
rect 24860 15020 24912 15026
rect 24492 14612 24544 14618
rect 24492 14554 24544 14560
rect 24504 14278 24532 14554
rect 24688 14346 24716 15014
rect 24860 14962 24912 14968
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 24780 14550 24808 14826
rect 24768 14544 24820 14550
rect 24768 14486 24820 14492
rect 24676 14340 24728 14346
rect 24676 14282 24728 14288
rect 24492 14272 24544 14278
rect 24492 14214 24544 14220
rect 24492 14000 24544 14006
rect 24492 13942 24544 13948
rect 24504 13394 24532 13942
rect 24688 13734 24716 14282
rect 24584 13728 24636 13734
rect 24584 13670 24636 13676
rect 24676 13728 24728 13734
rect 24676 13670 24728 13676
rect 24492 13388 24544 13394
rect 24492 13330 24544 13336
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24504 11694 24532 12718
rect 24596 12374 24624 13670
rect 24780 13546 24808 14486
rect 24872 14346 24900 14962
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25056 14482 25084 14758
rect 25044 14476 25096 14482
rect 25044 14418 25096 14424
rect 24860 14340 24912 14346
rect 24860 14282 24912 14288
rect 24780 13518 24900 13546
rect 24768 13388 24820 13394
rect 24768 13330 24820 13336
rect 24676 13320 24728 13326
rect 24676 13262 24728 13268
rect 24688 12646 24716 13262
rect 24780 12986 24808 13330
rect 24768 12980 24820 12986
rect 24768 12922 24820 12928
rect 24872 12866 24900 13518
rect 24952 13184 25004 13190
rect 24952 13126 25004 13132
rect 24780 12838 24900 12866
rect 24676 12640 24728 12646
rect 24676 12582 24728 12588
rect 24688 12442 24716 12582
rect 24676 12436 24728 12442
rect 24676 12378 24728 12384
rect 24584 12368 24636 12374
rect 24584 12310 24636 12316
rect 24780 11778 24808 12838
rect 24964 12238 24992 13126
rect 25056 12374 25084 14418
rect 25044 12368 25096 12374
rect 25044 12310 25096 12316
rect 24952 12232 25004 12238
rect 24952 12174 25004 12180
rect 24860 12164 24912 12170
rect 24860 12106 24912 12112
rect 24596 11750 24808 11778
rect 24492 11688 24544 11694
rect 24492 11630 24544 11636
rect 24400 11076 24452 11082
rect 24400 11018 24452 11024
rect 24412 10130 24440 11018
rect 24596 10538 24624 11750
rect 24676 11688 24728 11694
rect 24676 11630 24728 11636
rect 24584 10532 24636 10538
rect 24584 10474 24636 10480
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24412 9722 24440 10066
rect 24596 9926 24624 10474
rect 24688 10198 24716 11630
rect 24872 11626 24900 12106
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 24860 11620 24912 11626
rect 24860 11562 24912 11568
rect 24676 10192 24728 10198
rect 24676 10134 24728 10140
rect 24584 9920 24636 9926
rect 24584 9862 24636 9868
rect 24400 9716 24452 9722
rect 24400 9658 24452 9664
rect 24492 7744 24544 7750
rect 24492 7686 24544 7692
rect 24504 6730 24532 7686
rect 25056 7206 25084 11698
rect 25148 9994 25176 16730
rect 25136 9988 25188 9994
rect 25136 9930 25188 9936
rect 25240 7546 25268 21966
rect 25332 18612 25360 22510
rect 25424 22114 25452 28966
rect 25516 28762 25544 30654
rect 25596 30592 25648 30598
rect 25596 30534 25648 30540
rect 25608 29578 25636 30534
rect 25780 30184 25832 30190
rect 25780 30126 25832 30132
rect 25792 29782 25820 30126
rect 25780 29776 25832 29782
rect 25780 29718 25832 29724
rect 25596 29572 25648 29578
rect 25596 29514 25648 29520
rect 25780 29096 25832 29102
rect 25780 29038 25832 29044
rect 25504 28756 25556 28762
rect 25504 28698 25556 28704
rect 25516 28218 25544 28698
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25504 28212 25556 28218
rect 25504 28154 25556 28160
rect 25504 25832 25556 25838
rect 25504 25774 25556 25780
rect 25516 22234 25544 25774
rect 25504 22228 25556 22234
rect 25504 22170 25556 22176
rect 25424 22086 25544 22114
rect 25412 21956 25464 21962
rect 25412 21898 25464 21904
rect 25424 21486 25452 21898
rect 25412 21480 25464 21486
rect 25412 21422 25464 21428
rect 25412 19372 25464 19378
rect 25412 19314 25464 19320
rect 25516 19334 25544 22086
rect 25608 22094 25636 28562
rect 25688 28416 25740 28422
rect 25688 28358 25740 28364
rect 25700 28082 25728 28358
rect 25688 28076 25740 28082
rect 25688 28018 25740 28024
rect 25688 27668 25740 27674
rect 25688 27610 25740 27616
rect 25700 27418 25728 27610
rect 25792 27538 25820 29038
rect 25884 28966 25912 30806
rect 26056 30728 26108 30734
rect 26056 30670 26108 30676
rect 26068 30394 26096 30670
rect 26056 30388 26108 30394
rect 26056 30330 26108 30336
rect 25872 28960 25924 28966
rect 25872 28902 25924 28908
rect 25872 28688 25924 28694
rect 25872 28630 25924 28636
rect 25884 28082 25912 28630
rect 25872 28076 25924 28082
rect 25872 28018 25924 28024
rect 26056 28008 26108 28014
rect 26056 27950 26108 27956
rect 25780 27532 25832 27538
rect 25780 27474 25832 27480
rect 25700 27390 25820 27418
rect 25688 26308 25740 26314
rect 25688 26250 25740 26256
rect 25700 24818 25728 26250
rect 25688 24812 25740 24818
rect 25688 24754 25740 24760
rect 25792 24698 25820 27390
rect 26068 26790 26096 27950
rect 26056 26784 26108 26790
rect 26056 26726 26108 26732
rect 25872 26512 25924 26518
rect 25872 26454 25924 26460
rect 25884 24818 25912 26454
rect 26068 26450 26096 26726
rect 26252 26450 26280 31350
rect 26344 30818 26372 31826
rect 26436 31414 26464 45766
rect 26424 31408 26476 31414
rect 26424 31350 26476 31356
rect 26344 30790 26464 30818
rect 26332 30728 26384 30734
rect 26332 30670 26384 30676
rect 26344 30326 26372 30670
rect 26436 30666 26464 30790
rect 26424 30660 26476 30666
rect 26424 30602 26476 30608
rect 26332 30320 26384 30326
rect 26332 30262 26384 30268
rect 26344 29646 26372 30262
rect 26332 29640 26384 29646
rect 26332 29582 26384 29588
rect 26344 26994 26372 29582
rect 26332 26988 26384 26994
rect 26332 26930 26384 26936
rect 26424 26920 26476 26926
rect 26424 26862 26476 26868
rect 26056 26444 26108 26450
rect 26056 26386 26108 26392
rect 26240 26444 26292 26450
rect 26240 26386 26292 26392
rect 26148 26376 26200 26382
rect 26148 26318 26200 26324
rect 26056 25968 26108 25974
rect 26056 25910 26108 25916
rect 25872 24812 25924 24818
rect 25872 24754 25924 24760
rect 25700 24670 25820 24698
rect 25700 23322 25728 24670
rect 25872 24608 25924 24614
rect 25870 24576 25872 24585
rect 25924 24576 25926 24585
rect 25870 24511 25926 24520
rect 25872 24132 25924 24138
rect 25872 24074 25924 24080
rect 25884 23866 25912 24074
rect 25872 23860 25924 23866
rect 25872 23802 25924 23808
rect 25872 23724 25924 23730
rect 25872 23666 25924 23672
rect 25780 23656 25832 23662
rect 25780 23598 25832 23604
rect 25688 23316 25740 23322
rect 25688 23258 25740 23264
rect 25792 22438 25820 23598
rect 25780 22432 25832 22438
rect 25780 22374 25832 22380
rect 25608 22066 25728 22094
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25608 19854 25636 21966
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25700 19417 25728 22066
rect 25792 21554 25820 22374
rect 25780 21548 25832 21554
rect 25780 21490 25832 21496
rect 25780 19984 25832 19990
rect 25780 19926 25832 19932
rect 25686 19408 25742 19417
rect 25686 19343 25742 19352
rect 25424 18970 25452 19314
rect 25516 19306 25636 19334
rect 25412 18964 25464 18970
rect 25412 18906 25464 18912
rect 25412 18760 25464 18766
rect 25464 18708 25544 18714
rect 25412 18702 25544 18708
rect 25424 18686 25544 18702
rect 25332 18584 25452 18612
rect 25318 18320 25374 18329
rect 25318 18255 25320 18264
rect 25372 18255 25374 18264
rect 25320 18226 25372 18232
rect 25320 18080 25372 18086
rect 25320 18022 25372 18028
rect 25332 17610 25360 18022
rect 25320 17604 25372 17610
rect 25320 17546 25372 17552
rect 25332 16590 25360 17546
rect 25320 16584 25372 16590
rect 25320 16526 25372 16532
rect 25320 16040 25372 16046
rect 25320 15982 25372 15988
rect 25332 15570 25360 15982
rect 25320 15564 25372 15570
rect 25320 15506 25372 15512
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25332 12850 25360 13262
rect 25320 12844 25372 12850
rect 25320 12786 25372 12792
rect 25332 12306 25360 12786
rect 25320 12300 25372 12306
rect 25320 12242 25372 12248
rect 25332 11898 25360 12242
rect 25320 11892 25372 11898
rect 25320 11834 25372 11840
rect 25228 7540 25280 7546
rect 25228 7482 25280 7488
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 24964 6798 24992 7142
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24492 6724 24544 6730
rect 24492 6666 24544 6672
rect 25056 6390 25084 7142
rect 25044 6384 25096 6390
rect 25044 6326 25096 6332
rect 25424 5914 25452 18584
rect 25516 15978 25544 18686
rect 25608 18306 25636 19306
rect 25792 18698 25820 19926
rect 25884 18902 25912 23666
rect 25964 23316 26016 23322
rect 25964 23258 26016 23264
rect 25872 18896 25924 18902
rect 25872 18838 25924 18844
rect 25780 18692 25832 18698
rect 25780 18634 25832 18640
rect 25792 18426 25820 18634
rect 25780 18420 25832 18426
rect 25780 18362 25832 18368
rect 25872 18352 25924 18358
rect 25608 18278 25820 18306
rect 25872 18294 25924 18300
rect 25686 18184 25742 18193
rect 25686 18119 25742 18128
rect 25700 16454 25728 18119
rect 25688 16448 25740 16454
rect 25688 16390 25740 16396
rect 25504 15972 25556 15978
rect 25504 15914 25556 15920
rect 25596 15904 25648 15910
rect 25596 15846 25648 15852
rect 25608 15706 25636 15846
rect 25596 15700 25648 15706
rect 25596 15642 25648 15648
rect 25608 15586 25636 15642
rect 25608 15558 25728 15586
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25516 15162 25544 15438
rect 25504 15156 25556 15162
rect 25504 15098 25556 15104
rect 25504 13388 25556 13394
rect 25504 13330 25556 13336
rect 25516 11626 25544 13330
rect 25596 12912 25648 12918
rect 25596 12854 25648 12860
rect 25608 12102 25636 12854
rect 25596 12096 25648 12102
rect 25596 12038 25648 12044
rect 25596 11688 25648 11694
rect 25596 11630 25648 11636
rect 25504 11620 25556 11626
rect 25504 11562 25556 11568
rect 25608 11354 25636 11630
rect 25700 11354 25728 15558
rect 25792 11762 25820 18278
rect 25884 17678 25912 18294
rect 25872 17672 25924 17678
rect 25872 17614 25924 17620
rect 25872 17128 25924 17134
rect 25872 17070 25924 17076
rect 25780 11756 25832 11762
rect 25780 11698 25832 11704
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25688 11348 25740 11354
rect 25688 11290 25740 11296
rect 25780 9920 25832 9926
rect 25780 9862 25832 9868
rect 25792 9586 25820 9862
rect 25780 9580 25832 9586
rect 25780 9522 25832 9528
rect 25792 9178 25820 9522
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25884 7562 25912 17070
rect 25976 16794 26004 23258
rect 26068 19904 26096 25910
rect 26160 25906 26188 26318
rect 26148 25900 26200 25906
rect 26148 25842 26200 25848
rect 26160 25498 26188 25842
rect 26148 25492 26200 25498
rect 26148 25434 26200 25440
rect 26160 25294 26188 25434
rect 26148 25288 26200 25294
rect 26148 25230 26200 25236
rect 26252 25226 26280 26386
rect 26436 26314 26464 26862
rect 26424 26308 26476 26314
rect 26424 26250 26476 26256
rect 26240 25220 26292 25226
rect 26240 25162 26292 25168
rect 26436 24732 26464 26250
rect 26344 24704 26464 24732
rect 26238 23624 26294 23633
rect 26238 23559 26294 23568
rect 26252 23526 26280 23559
rect 26240 23520 26292 23526
rect 26240 23462 26292 23468
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22710 26280 22918
rect 26240 22704 26292 22710
rect 26240 22646 26292 22652
rect 26344 22094 26372 24704
rect 26424 24608 26476 24614
rect 26424 24550 26476 24556
rect 26252 22066 26372 22094
rect 26252 21690 26280 22066
rect 26240 21684 26292 21690
rect 26240 21626 26292 21632
rect 26148 21616 26200 21622
rect 26148 21558 26200 21564
rect 26160 20874 26188 21558
rect 26240 20936 26292 20942
rect 26240 20878 26292 20884
rect 26148 20868 26200 20874
rect 26148 20810 26200 20816
rect 26252 20505 26280 20878
rect 26238 20496 26294 20505
rect 26238 20431 26294 20440
rect 26068 19876 26188 19904
rect 26056 19780 26108 19786
rect 26056 19722 26108 19728
rect 26068 19514 26096 19722
rect 26056 19508 26108 19514
rect 26056 19450 26108 19456
rect 26160 19394 26188 19876
rect 26068 19366 26188 19394
rect 26068 18329 26096 19366
rect 26436 19310 26464 24550
rect 26424 19304 26476 19310
rect 26330 19272 26386 19281
rect 26424 19246 26476 19252
rect 26330 19207 26386 19216
rect 26240 18896 26292 18902
rect 26240 18838 26292 18844
rect 26148 18760 26200 18766
rect 26148 18702 26200 18708
rect 26054 18320 26110 18329
rect 26054 18255 26110 18264
rect 26056 18216 26108 18222
rect 26056 18158 26108 18164
rect 26068 17202 26096 18158
rect 26160 17882 26188 18702
rect 26252 18290 26280 18838
rect 26240 18284 26292 18290
rect 26240 18226 26292 18232
rect 26148 17876 26200 17882
rect 26148 17818 26200 17824
rect 26344 17338 26372 19207
rect 26436 18970 26464 19246
rect 26424 18964 26476 18970
rect 26424 18906 26476 18912
rect 26332 17332 26384 17338
rect 26160 17292 26332 17320
rect 26056 17196 26108 17202
rect 26056 17138 26108 17144
rect 25964 16788 26016 16794
rect 25964 16730 26016 16736
rect 26056 16516 26108 16522
rect 26056 16458 26108 16464
rect 26068 15570 26096 16458
rect 26160 16153 26188 17292
rect 26332 17274 26384 17280
rect 26436 16658 26464 18906
rect 26424 16652 26476 16658
rect 26424 16594 26476 16600
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26146 16144 26202 16153
rect 26146 16079 26202 16088
rect 26056 15564 26108 15570
rect 26056 15506 26108 15512
rect 26056 15360 26108 15366
rect 26056 15302 26108 15308
rect 25964 13456 26016 13462
rect 25964 13398 26016 13404
rect 25976 9654 26004 13398
rect 26068 12832 26096 15302
rect 26160 15026 26188 16079
rect 26332 15904 26384 15910
rect 26332 15846 26384 15852
rect 26344 15434 26372 15846
rect 26332 15428 26384 15434
rect 26332 15370 26384 15376
rect 26148 15020 26200 15026
rect 26148 14962 26200 14968
rect 26240 14952 26292 14958
rect 26240 14894 26292 14900
rect 26148 14272 26200 14278
rect 26148 14214 26200 14220
rect 26160 14006 26188 14214
rect 26148 14000 26200 14006
rect 26148 13942 26200 13948
rect 26252 13462 26280 14894
rect 26436 14618 26464 16390
rect 26528 15994 26556 47670
rect 27160 47660 27212 47666
rect 27160 47602 27212 47608
rect 26700 43784 26752 43790
rect 26700 43726 26752 43732
rect 26608 40180 26660 40186
rect 26608 40122 26660 40128
rect 26620 39409 26648 40122
rect 26606 39400 26662 39409
rect 26606 39335 26662 39344
rect 26620 34746 26648 39335
rect 26608 34740 26660 34746
rect 26608 34682 26660 34688
rect 26608 34604 26660 34610
rect 26608 34546 26660 34552
rect 26620 34066 26648 34546
rect 26608 34060 26660 34066
rect 26608 34002 26660 34008
rect 26712 27010 26740 43726
rect 27068 37188 27120 37194
rect 27068 37130 27120 37136
rect 26976 36780 27028 36786
rect 26976 36722 27028 36728
rect 26792 36304 26844 36310
rect 26792 36246 26844 36252
rect 26804 35154 26832 36246
rect 26884 36100 26936 36106
rect 26884 36042 26936 36048
rect 26792 35148 26844 35154
rect 26792 35090 26844 35096
rect 26792 32224 26844 32230
rect 26792 32166 26844 32172
rect 26804 31822 26832 32166
rect 26792 31816 26844 31822
rect 26792 31758 26844 31764
rect 26804 31482 26832 31758
rect 26792 31476 26844 31482
rect 26792 31418 26844 31424
rect 26792 30932 26844 30938
rect 26792 30874 26844 30880
rect 26804 27538 26832 30874
rect 26792 27532 26844 27538
rect 26792 27474 26844 27480
rect 26712 26982 26832 27010
rect 26700 26784 26752 26790
rect 26700 26726 26752 26732
rect 26606 24304 26662 24313
rect 26606 24239 26662 24248
rect 26620 23798 26648 24239
rect 26608 23792 26660 23798
rect 26608 23734 26660 23740
rect 26608 20324 26660 20330
rect 26608 20266 26660 20272
rect 26620 19922 26648 20266
rect 26608 19916 26660 19922
rect 26608 19858 26660 19864
rect 26608 19168 26660 19174
rect 26608 19110 26660 19116
rect 26620 18698 26648 19110
rect 26608 18692 26660 18698
rect 26608 18634 26660 18640
rect 26528 15966 26648 15994
rect 26516 15360 26568 15366
rect 26516 15302 26568 15308
rect 26528 15026 26556 15302
rect 26516 15020 26568 15026
rect 26516 14962 26568 14968
rect 26424 14612 26476 14618
rect 26424 14554 26476 14560
rect 26436 13870 26464 14554
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26332 13796 26384 13802
rect 26332 13738 26384 13744
rect 26240 13456 26292 13462
rect 26240 13398 26292 13404
rect 26240 12844 26292 12850
rect 26068 12804 26240 12832
rect 26240 12786 26292 12792
rect 26252 12753 26280 12786
rect 26344 12782 26372 13738
rect 26332 12776 26384 12782
rect 26238 12744 26294 12753
rect 26148 12708 26200 12714
rect 26332 12718 26384 12724
rect 26238 12679 26294 12688
rect 26148 12650 26200 12656
rect 26160 12102 26188 12650
rect 26424 12640 26476 12646
rect 26424 12582 26476 12588
rect 26436 12170 26464 12582
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26056 12096 26108 12102
rect 26056 12038 26108 12044
rect 26148 12096 26200 12102
rect 26148 12038 26200 12044
rect 26068 11898 26096 12038
rect 26056 11892 26108 11898
rect 26056 11834 26108 11840
rect 26160 11694 26188 12038
rect 26148 11688 26200 11694
rect 26148 11630 26200 11636
rect 26332 11688 26384 11694
rect 26332 11630 26384 11636
rect 26240 11348 26292 11354
rect 26240 11290 26292 11296
rect 26252 10674 26280 11290
rect 26344 11218 26372 11630
rect 26332 11212 26384 11218
rect 26332 11154 26384 11160
rect 26240 10668 26292 10674
rect 26240 10610 26292 10616
rect 26252 10266 26280 10610
rect 26332 10600 26384 10606
rect 26384 10548 26464 10554
rect 26332 10542 26464 10548
rect 26344 10526 26464 10542
rect 26332 10464 26384 10470
rect 26332 10406 26384 10412
rect 26240 10260 26292 10266
rect 26240 10202 26292 10208
rect 26056 9988 26108 9994
rect 26056 9930 26108 9936
rect 25964 9648 26016 9654
rect 25964 9590 26016 9596
rect 25976 9042 26004 9590
rect 26068 9518 26096 9930
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 26344 9450 26372 10406
rect 26436 10266 26464 10526
rect 26516 10464 26568 10470
rect 26516 10406 26568 10412
rect 26424 10260 26476 10266
rect 26424 10202 26476 10208
rect 26528 10130 26556 10406
rect 26516 10124 26568 10130
rect 26516 10066 26568 10072
rect 26424 9920 26476 9926
rect 26424 9862 26476 9868
rect 26436 9586 26464 9862
rect 26528 9654 26556 10066
rect 26516 9648 26568 9654
rect 26516 9590 26568 9596
rect 26424 9580 26476 9586
rect 26424 9522 26476 9528
rect 26332 9444 26384 9450
rect 26332 9386 26384 9392
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 25964 9036 26016 9042
rect 25964 8978 26016 8984
rect 25792 7534 25912 7562
rect 25412 5908 25464 5914
rect 25412 5850 25464 5856
rect 24398 4040 24454 4049
rect 24398 3975 24400 3984
rect 24452 3975 24454 3984
rect 24400 3946 24452 3952
rect 25688 3936 25740 3942
rect 25688 3878 25740 3884
rect 25700 3602 25728 3878
rect 25504 3596 25556 3602
rect 25504 3538 25556 3544
rect 25688 3596 25740 3602
rect 25688 3538 25740 3544
rect 25516 3126 25544 3538
rect 25504 3120 25556 3126
rect 25504 3062 25556 3068
rect 24136 2746 24256 2774
rect 24136 2582 24164 2746
rect 24124 2576 24176 2582
rect 24124 2518 24176 2524
rect 23940 2508 23992 2514
rect 23940 2450 23992 2456
rect 24492 2440 24544 2446
rect 24492 2382 24544 2388
rect 25136 2440 25188 2446
rect 25136 2382 25188 2388
rect 24504 800 24532 2382
rect 25148 800 25176 2382
rect 25792 2378 25820 7534
rect 25976 7342 26004 8978
rect 26252 8974 26280 9318
rect 26240 8968 26292 8974
rect 26240 8910 26292 8916
rect 26436 8430 26464 9522
rect 26424 8424 26476 8430
rect 26424 8366 26476 8372
rect 26620 7970 26648 15966
rect 26436 7942 26648 7970
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 25976 6798 26004 7278
rect 25964 6792 26016 6798
rect 25964 6734 26016 6740
rect 25872 5704 25924 5710
rect 25872 5646 25924 5652
rect 25884 2582 25912 5646
rect 26436 4078 26464 7942
rect 26712 7834 26740 26726
rect 26804 26058 26832 26982
rect 26896 26790 26924 36042
rect 26988 34134 27016 36722
rect 27080 36582 27108 37130
rect 27068 36576 27120 36582
rect 27068 36518 27120 36524
rect 27172 35986 27200 47602
rect 27344 40112 27396 40118
rect 27344 40054 27396 40060
rect 27356 39030 27384 40054
rect 27528 39976 27580 39982
rect 27528 39918 27580 39924
rect 27344 39024 27396 39030
rect 27344 38966 27396 38972
rect 27356 38842 27384 38966
rect 27540 38894 27568 39918
rect 27264 38814 27384 38842
rect 27528 38888 27580 38894
rect 27528 38830 27580 38836
rect 27264 37670 27292 38814
rect 27344 38752 27396 38758
rect 27344 38694 27396 38700
rect 27356 38350 27384 38694
rect 27344 38344 27396 38350
rect 27344 38286 27396 38292
rect 27252 37664 27304 37670
rect 27252 37606 27304 37612
rect 27528 36168 27580 36174
rect 27526 36136 27528 36145
rect 27580 36136 27582 36145
rect 27526 36071 27582 36080
rect 27080 35958 27200 35986
rect 26976 34128 27028 34134
rect 26976 34070 27028 34076
rect 26988 32910 27016 34070
rect 26976 32904 27028 32910
rect 26976 32846 27028 32852
rect 26976 31136 27028 31142
rect 26976 31078 27028 31084
rect 26988 30734 27016 31078
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 27080 28762 27108 35958
rect 27436 35692 27488 35698
rect 27436 35634 27488 35640
rect 27344 35556 27396 35562
rect 27344 35498 27396 35504
rect 27252 35488 27304 35494
rect 27252 35430 27304 35436
rect 27264 35086 27292 35430
rect 27252 35080 27304 35086
rect 27252 35022 27304 35028
rect 27356 34678 27384 35498
rect 27448 35290 27476 35634
rect 27436 35284 27488 35290
rect 27436 35226 27488 35232
rect 27540 35086 27568 36071
rect 27618 35592 27674 35601
rect 27618 35527 27674 35536
rect 27632 35290 27660 35527
rect 27620 35284 27672 35290
rect 27620 35226 27672 35232
rect 27528 35080 27580 35086
rect 27528 35022 27580 35028
rect 27528 34944 27580 34950
rect 27528 34886 27580 34892
rect 27344 34672 27396 34678
rect 27344 34614 27396 34620
rect 27160 33584 27212 33590
rect 27158 33552 27160 33561
rect 27212 33552 27214 33561
rect 27158 33487 27214 33496
rect 27160 33312 27212 33318
rect 27160 33254 27212 33260
rect 27172 33046 27200 33254
rect 27160 33040 27212 33046
rect 27160 32982 27212 32988
rect 27344 32360 27396 32366
rect 27344 32302 27396 32308
rect 27160 31884 27212 31890
rect 27160 31826 27212 31832
rect 27172 31686 27200 31826
rect 27160 31680 27212 31686
rect 27160 31622 27212 31628
rect 27172 31142 27200 31622
rect 27160 31136 27212 31142
rect 27160 31078 27212 31084
rect 27356 29714 27384 32302
rect 27344 29708 27396 29714
rect 27344 29650 27396 29656
rect 27252 29640 27304 29646
rect 27252 29582 27304 29588
rect 27068 28756 27120 28762
rect 27068 28698 27120 28704
rect 27264 28694 27292 29582
rect 27252 28688 27304 28694
rect 27252 28630 27304 28636
rect 27434 28112 27490 28121
rect 27434 28047 27436 28056
rect 27488 28047 27490 28056
rect 27436 28018 27488 28024
rect 27344 27872 27396 27878
rect 27344 27814 27396 27820
rect 27356 27470 27384 27814
rect 27252 27464 27304 27470
rect 27252 27406 27304 27412
rect 27344 27464 27396 27470
rect 27344 27406 27396 27412
rect 27264 26994 27292 27406
rect 27434 27024 27490 27033
rect 27252 26988 27304 26994
rect 27434 26959 27436 26968
rect 27252 26930 27304 26936
rect 27488 26959 27490 26968
rect 27436 26930 27488 26936
rect 26884 26784 26936 26790
rect 26884 26726 26936 26732
rect 27252 26784 27304 26790
rect 27252 26726 27304 26732
rect 27264 26382 27292 26726
rect 27252 26376 27304 26382
rect 27252 26318 27304 26324
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 26804 26030 27016 26058
rect 26988 25974 27016 26030
rect 26976 25968 27028 25974
rect 26976 25910 27028 25916
rect 27160 25696 27212 25702
rect 27160 25638 27212 25644
rect 27172 25430 27200 25638
rect 27160 25424 27212 25430
rect 27160 25366 27212 25372
rect 26976 25152 27028 25158
rect 26976 25094 27028 25100
rect 26988 24954 27016 25094
rect 27158 24984 27214 24993
rect 26976 24948 27028 24954
rect 27158 24919 27214 24928
rect 26976 24890 27028 24896
rect 27172 24750 27200 24919
rect 27356 24818 27384 26182
rect 27436 25220 27488 25226
rect 27436 25162 27488 25168
rect 27344 24812 27396 24818
rect 27344 24754 27396 24760
rect 27160 24744 27212 24750
rect 27160 24686 27212 24692
rect 27160 24064 27212 24070
rect 27160 24006 27212 24012
rect 27172 23730 27200 24006
rect 26792 23724 26844 23730
rect 26792 23666 26844 23672
rect 26976 23724 27028 23730
rect 26976 23666 27028 23672
rect 27160 23724 27212 23730
rect 27160 23666 27212 23672
rect 26804 23594 26832 23666
rect 26792 23588 26844 23594
rect 26792 23530 26844 23536
rect 26804 19990 26832 23530
rect 26988 23050 27016 23666
rect 26976 23044 27028 23050
rect 26976 22986 27028 22992
rect 27252 23044 27304 23050
rect 27252 22986 27304 22992
rect 26884 22704 26936 22710
rect 26884 22646 26936 22652
rect 26792 19984 26844 19990
rect 26792 19926 26844 19932
rect 26792 19712 26844 19718
rect 26792 19654 26844 19660
rect 26804 14770 26832 19654
rect 26896 18034 26924 22646
rect 26988 21622 27016 22986
rect 27264 22642 27292 22986
rect 27252 22636 27304 22642
rect 27252 22578 27304 22584
rect 27448 22094 27476 25162
rect 27356 22066 27476 22094
rect 27160 21888 27212 21894
rect 27160 21830 27212 21836
rect 26976 21616 27028 21622
rect 26976 21558 27028 21564
rect 27172 21554 27200 21830
rect 27160 21548 27212 21554
rect 27160 21490 27212 21496
rect 27172 21010 27200 21490
rect 27160 21004 27212 21010
rect 27160 20946 27212 20952
rect 26896 18006 27016 18034
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 26896 15366 26924 17818
rect 26988 16590 27016 18006
rect 27160 16652 27212 16658
rect 27160 16594 27212 16600
rect 26976 16584 27028 16590
rect 26976 16526 27028 16532
rect 27172 16114 27200 16594
rect 27252 16584 27304 16590
rect 27252 16526 27304 16532
rect 26976 16108 27028 16114
rect 26976 16050 27028 16056
rect 27160 16108 27212 16114
rect 27160 16050 27212 16056
rect 26988 15706 27016 16050
rect 26976 15700 27028 15706
rect 26976 15642 27028 15648
rect 27172 15502 27200 16050
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26884 15360 26936 15366
rect 26884 15302 26936 15308
rect 26896 14890 26924 15302
rect 26884 14884 26936 14890
rect 26884 14826 26936 14832
rect 26804 14742 26924 14770
rect 26896 14006 26924 14742
rect 26884 14000 26936 14006
rect 26884 13942 26936 13948
rect 26896 12646 26924 13942
rect 27264 13938 27292 16526
rect 27252 13932 27304 13938
rect 27252 13874 27304 13880
rect 27264 13530 27292 13874
rect 27252 13524 27304 13530
rect 27252 13466 27304 13472
rect 27160 13388 27212 13394
rect 27160 13330 27212 13336
rect 27172 12986 27200 13330
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27160 12980 27212 12986
rect 27160 12922 27212 12928
rect 27264 12850 27292 13126
rect 27252 12844 27304 12850
rect 27252 12786 27304 12792
rect 27250 12744 27306 12753
rect 27250 12679 27306 12688
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 27172 12322 27200 12582
rect 27264 12374 27292 12679
rect 26988 12294 27200 12322
rect 27252 12368 27304 12374
rect 27252 12310 27304 12316
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26804 10033 26832 11834
rect 26790 10024 26846 10033
rect 26790 9959 26846 9968
rect 26528 7806 26740 7834
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26424 3596 26476 3602
rect 26424 3538 26476 3544
rect 26148 3460 26200 3466
rect 26148 3402 26200 3408
rect 26160 2854 26188 3402
rect 26148 2848 26200 2854
rect 26148 2790 26200 2796
rect 25872 2576 25924 2582
rect 25872 2518 25924 2524
rect 25780 2372 25832 2378
rect 25780 2314 25832 2320
rect 26436 800 26464 3538
rect 26528 1902 26556 7806
rect 26608 7744 26660 7750
rect 26608 7686 26660 7692
rect 26620 7478 26648 7686
rect 26608 7472 26660 7478
rect 26608 7414 26660 7420
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26712 6866 26740 7142
rect 26700 6860 26752 6866
rect 26700 6802 26752 6808
rect 26804 5574 26832 9959
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26896 7886 26924 8842
rect 26884 7880 26936 7886
rect 26884 7822 26936 7828
rect 26896 7002 26924 7822
rect 26988 7750 27016 12294
rect 27356 11898 27384 22066
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27448 17134 27476 17614
rect 27436 17128 27488 17134
rect 27436 17070 27488 17076
rect 27448 15094 27476 17070
rect 27436 15088 27488 15094
rect 27436 15030 27488 15036
rect 27540 15026 27568 34886
rect 27724 29594 27752 49098
rect 27816 48686 27844 51326
rect 28354 51326 28488 51354
rect 28354 51200 28410 51326
rect 27988 49224 28040 49230
rect 27988 49166 28040 49172
rect 27804 48680 27856 48686
rect 27804 48622 27856 48628
rect 28000 47666 28028 49166
rect 27988 47660 28040 47666
rect 27988 47602 28040 47608
rect 28460 47598 28488 51326
rect 28998 51200 29054 52000
rect 29642 51354 29698 52000
rect 29642 51326 29868 51354
rect 29642 51200 29698 51326
rect 29012 49230 29040 51200
rect 29000 49224 29052 49230
rect 29000 49166 29052 49172
rect 29840 48686 29868 51326
rect 30930 51200 30986 52000
rect 31574 51200 31630 52000
rect 32218 51200 32274 52000
rect 32862 51354 32918 52000
rect 32862 51326 33088 51354
rect 32862 51200 32918 51326
rect 29920 49360 29972 49366
rect 29920 49302 29972 49308
rect 29276 48680 29328 48686
rect 29276 48622 29328 48628
rect 29552 48680 29604 48686
rect 29552 48622 29604 48628
rect 29828 48680 29880 48686
rect 29828 48622 29880 48628
rect 28172 47592 28224 47598
rect 28172 47534 28224 47540
rect 28448 47592 28500 47598
rect 28448 47534 28500 47540
rect 28184 47258 28212 47534
rect 28172 47252 28224 47258
rect 28172 47194 28224 47200
rect 28264 47048 28316 47054
rect 28264 46990 28316 46996
rect 28276 45558 28304 46990
rect 28264 45552 28316 45558
rect 28264 45494 28316 45500
rect 28080 40044 28132 40050
rect 28080 39986 28132 39992
rect 28092 39574 28120 39986
rect 28080 39568 28132 39574
rect 28080 39510 28132 39516
rect 27804 39296 27856 39302
rect 27804 39238 27856 39244
rect 27816 39098 27844 39238
rect 27804 39092 27856 39098
rect 27804 39034 27856 39040
rect 27804 38956 27856 38962
rect 27804 38898 27856 38904
rect 27816 38554 27844 38898
rect 27804 38548 27856 38554
rect 27804 38490 27856 38496
rect 27816 37806 27844 38490
rect 28092 38418 28120 39510
rect 28080 38412 28132 38418
rect 28080 38354 28132 38360
rect 27804 37800 27856 37806
rect 27804 37742 27856 37748
rect 27804 37392 27856 37398
rect 27804 37334 27856 37340
rect 27816 36786 27844 37334
rect 27804 36780 27856 36786
rect 27804 36722 27856 36728
rect 27896 36780 27948 36786
rect 27896 36722 27948 36728
rect 27816 35766 27844 36722
rect 27908 36378 27936 36722
rect 27896 36372 27948 36378
rect 27896 36314 27948 36320
rect 27804 35760 27856 35766
rect 27804 35702 27856 35708
rect 27988 35012 28040 35018
rect 27988 34954 28040 34960
rect 27804 34468 27856 34474
rect 27804 34410 27856 34416
rect 27816 29646 27844 34410
rect 28000 33998 28028 34954
rect 28092 34610 28120 38354
rect 28172 36304 28224 36310
rect 28172 36246 28224 36252
rect 28080 34604 28132 34610
rect 28080 34546 28132 34552
rect 28184 34474 28212 36246
rect 28172 34468 28224 34474
rect 28172 34410 28224 34416
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 28092 34202 28120 34342
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 27988 33992 28040 33998
rect 27988 33934 28040 33940
rect 27896 32836 27948 32842
rect 27896 32778 27948 32784
rect 27908 32502 27936 32778
rect 27896 32496 27948 32502
rect 27896 32438 27948 32444
rect 27908 31414 27936 32438
rect 27896 31408 27948 31414
rect 27896 31350 27948 31356
rect 27632 29566 27752 29594
rect 27804 29640 27856 29646
rect 27804 29582 27856 29588
rect 27632 26790 27660 29566
rect 27712 29504 27764 29510
rect 27712 29446 27764 29452
rect 27724 28218 27752 29446
rect 27988 28484 28040 28490
rect 27988 28426 28040 28432
rect 27894 28384 27950 28393
rect 27894 28319 27950 28328
rect 27712 28212 27764 28218
rect 27712 28154 27764 28160
rect 27908 27946 27936 28319
rect 27896 27940 27948 27946
rect 27896 27882 27948 27888
rect 28000 27305 28028 28426
rect 28092 28121 28120 34138
rect 28172 29708 28224 29714
rect 28172 29650 28224 29656
rect 28184 28626 28212 29650
rect 28172 28620 28224 28626
rect 28172 28562 28224 28568
rect 28078 28112 28134 28121
rect 28078 28047 28134 28056
rect 27986 27296 28042 27305
rect 27986 27231 28042 27240
rect 28172 26988 28224 26994
rect 28172 26930 28224 26936
rect 27620 26784 27672 26790
rect 27620 26726 27672 26732
rect 28184 26042 28212 26930
rect 28172 26036 28224 26042
rect 28172 25978 28224 25984
rect 27988 25696 28040 25702
rect 27988 25638 28040 25644
rect 28000 25294 28028 25638
rect 27988 25288 28040 25294
rect 27988 25230 28040 25236
rect 28000 24818 28028 25230
rect 28276 25226 28304 45494
rect 29000 39976 29052 39982
rect 29000 39918 29052 39924
rect 28908 39840 28960 39846
rect 28908 39782 28960 39788
rect 28448 39500 28500 39506
rect 28448 39442 28500 39448
rect 28356 39296 28408 39302
rect 28356 39238 28408 39244
rect 28368 39030 28396 39238
rect 28356 39024 28408 39030
rect 28356 38966 28408 38972
rect 28460 38418 28488 39442
rect 28540 39432 28592 39438
rect 28540 39374 28592 39380
rect 28552 38962 28580 39374
rect 28920 39370 28948 39782
rect 29012 39438 29040 39918
rect 29000 39432 29052 39438
rect 29000 39374 29052 39380
rect 28908 39364 28960 39370
rect 28908 39306 28960 39312
rect 28816 39296 28868 39302
rect 28816 39238 28868 39244
rect 28540 38956 28592 38962
rect 28540 38898 28592 38904
rect 28552 38486 28580 38898
rect 28540 38480 28592 38486
rect 28540 38422 28592 38428
rect 28448 38412 28500 38418
rect 28448 38354 28500 38360
rect 28460 37738 28488 38354
rect 28448 37732 28500 37738
rect 28448 37674 28500 37680
rect 28552 37398 28580 38422
rect 28632 38344 28684 38350
rect 28632 38286 28684 38292
rect 28540 37392 28592 37398
rect 28540 37334 28592 37340
rect 28644 35034 28672 38286
rect 28644 35006 28764 35034
rect 28356 34400 28408 34406
rect 28356 34342 28408 34348
rect 28368 33998 28396 34342
rect 28356 33992 28408 33998
rect 28356 33934 28408 33940
rect 28368 33454 28396 33934
rect 28632 33924 28684 33930
rect 28632 33866 28684 33872
rect 28644 33658 28672 33866
rect 28632 33652 28684 33658
rect 28632 33594 28684 33600
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28368 32416 28396 33390
rect 28540 32904 28592 32910
rect 28540 32846 28592 32852
rect 28448 32428 28500 32434
rect 28368 32388 28448 32416
rect 28368 32026 28396 32388
rect 28448 32370 28500 32376
rect 28356 32020 28408 32026
rect 28356 31962 28408 31968
rect 28368 31754 28396 31962
rect 28356 31748 28408 31754
rect 28356 31690 28408 31696
rect 28448 29708 28500 29714
rect 28448 29650 28500 29656
rect 28460 29238 28488 29650
rect 28448 29232 28500 29238
rect 28448 29174 28500 29180
rect 28356 28416 28408 28422
rect 28356 28358 28408 28364
rect 28368 28082 28396 28358
rect 28356 28076 28408 28082
rect 28356 28018 28408 28024
rect 28448 26376 28500 26382
rect 28448 26318 28500 26324
rect 28460 26042 28488 26318
rect 28448 26036 28500 26042
rect 28448 25978 28500 25984
rect 28356 25968 28408 25974
rect 28408 25916 28488 25922
rect 28356 25910 28488 25916
rect 28368 25894 28488 25910
rect 28356 25492 28408 25498
rect 28356 25434 28408 25440
rect 28264 25220 28316 25226
rect 28264 25162 28316 25168
rect 27988 24812 28040 24818
rect 27988 24754 28040 24760
rect 27988 24608 28040 24614
rect 27988 24550 28040 24556
rect 27620 24200 27672 24206
rect 27620 24142 27672 24148
rect 28000 24188 28028 24550
rect 28368 24290 28396 25434
rect 28276 24262 28396 24290
rect 28172 24200 28224 24206
rect 28000 24160 28172 24188
rect 27632 22030 27660 24142
rect 27896 24132 27948 24138
rect 27896 24074 27948 24080
rect 27908 23866 27936 24074
rect 27896 23860 27948 23866
rect 27896 23802 27948 23808
rect 27804 23724 27856 23730
rect 27804 23666 27856 23672
rect 27620 22024 27672 22030
rect 27620 21966 27672 21972
rect 27816 21865 27844 23666
rect 28000 22094 28028 24160
rect 28172 24142 28224 24148
rect 28276 24018 28304 24262
rect 28356 24132 28408 24138
rect 28356 24074 28408 24080
rect 28184 23990 28304 24018
rect 28080 23656 28132 23662
rect 28080 23598 28132 23604
rect 28092 23254 28120 23598
rect 28080 23248 28132 23254
rect 28080 23190 28132 23196
rect 27908 22066 28028 22094
rect 27802 21856 27858 21865
rect 27724 21814 27802 21842
rect 27620 19848 27672 19854
rect 27620 19790 27672 19796
rect 27632 18290 27660 19790
rect 27620 18284 27672 18290
rect 27620 18226 27672 18232
rect 27724 18170 27752 21814
rect 27802 21791 27858 21800
rect 27804 19780 27856 19786
rect 27804 19722 27856 19728
rect 27816 18766 27844 19722
rect 27804 18760 27856 18766
rect 27804 18702 27856 18708
rect 27632 18142 27752 18170
rect 27632 17678 27660 18142
rect 27908 17898 27936 22066
rect 28092 21486 28120 23190
rect 28080 21480 28132 21486
rect 28080 21422 28132 21428
rect 27988 20800 28040 20806
rect 27988 20742 28040 20748
rect 28000 20534 28028 20742
rect 27988 20528 28040 20534
rect 27988 20470 28040 20476
rect 27988 18692 28040 18698
rect 27988 18634 28040 18640
rect 27724 17870 27936 17898
rect 27620 17672 27672 17678
rect 27620 17614 27672 17620
rect 27620 17264 27672 17270
rect 27620 17206 27672 17212
rect 27632 16590 27660 17206
rect 27620 16584 27672 16590
rect 27620 16526 27672 16532
rect 27618 15736 27674 15745
rect 27618 15671 27674 15680
rect 27528 15020 27580 15026
rect 27528 14962 27580 14968
rect 27436 14272 27488 14278
rect 27436 14214 27488 14220
rect 27448 14074 27476 14214
rect 27436 14068 27488 14074
rect 27436 14010 27488 14016
rect 27344 11892 27396 11898
rect 27344 11834 27396 11840
rect 27068 11756 27120 11762
rect 27068 11698 27120 11704
rect 27080 10538 27108 11698
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27160 11280 27212 11286
rect 27160 11222 27212 11228
rect 27172 10742 27200 11222
rect 27160 10736 27212 10742
rect 27160 10678 27212 10684
rect 27356 10674 27384 11290
rect 27344 10668 27396 10674
rect 27344 10610 27396 10616
rect 27068 10532 27120 10538
rect 27068 10474 27120 10480
rect 27344 10464 27396 10470
rect 27344 10406 27396 10412
rect 27356 9178 27384 10406
rect 27448 9330 27476 14010
rect 27632 12918 27660 15671
rect 27620 12912 27672 12918
rect 27620 12854 27672 12860
rect 27528 12232 27580 12238
rect 27528 12174 27580 12180
rect 27540 11286 27568 12174
rect 27632 11762 27660 12854
rect 27724 12434 27752 17870
rect 27896 17740 27948 17746
rect 27896 17682 27948 17688
rect 27804 16108 27856 16114
rect 27804 16050 27856 16056
rect 27816 15745 27844 16050
rect 27908 15978 27936 17682
rect 27896 15972 27948 15978
rect 27896 15914 27948 15920
rect 27802 15736 27858 15745
rect 27802 15671 27858 15680
rect 27896 15428 27948 15434
rect 27896 15370 27948 15376
rect 27908 15162 27936 15370
rect 27896 15156 27948 15162
rect 27896 15098 27948 15104
rect 27804 14340 27856 14346
rect 27804 14282 27856 14288
rect 27816 13326 27844 14282
rect 27908 13938 27936 15098
rect 28000 14414 28028 18634
rect 28184 18465 28212 23990
rect 28368 23866 28396 24074
rect 28356 23860 28408 23866
rect 28356 23802 28408 23808
rect 28356 23724 28408 23730
rect 28356 23666 28408 23672
rect 28368 23322 28396 23666
rect 28356 23316 28408 23322
rect 28356 23258 28408 23264
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28276 21690 28304 21898
rect 28264 21684 28316 21690
rect 28264 21626 28316 21632
rect 28170 18456 28226 18465
rect 28170 18391 28226 18400
rect 28080 17808 28132 17814
rect 28184 17785 28212 18391
rect 28264 18284 28316 18290
rect 28264 18226 28316 18232
rect 28080 17750 28132 17756
rect 28170 17776 28226 17785
rect 28092 16114 28120 17750
rect 28170 17711 28226 17720
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28184 17202 28212 17614
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28080 16108 28132 16114
rect 28080 16050 28132 16056
rect 28184 15638 28212 17138
rect 28276 16794 28304 18226
rect 28460 17921 28488 25894
rect 28446 17912 28502 17921
rect 28446 17847 28502 17856
rect 28448 17672 28500 17678
rect 28448 17614 28500 17620
rect 28356 17536 28408 17542
rect 28356 17478 28408 17484
rect 28264 16788 28316 16794
rect 28264 16730 28316 16736
rect 28368 16590 28396 17478
rect 28460 17134 28488 17614
rect 28448 17128 28500 17134
rect 28448 17070 28500 17076
rect 28356 16584 28408 16590
rect 28356 16526 28408 16532
rect 28354 16416 28410 16425
rect 28354 16351 28410 16360
rect 28172 15632 28224 15638
rect 28172 15574 28224 15580
rect 27988 14408 28040 14414
rect 27988 14350 28040 14356
rect 27896 13932 27948 13938
rect 27896 13874 27948 13880
rect 27908 13326 27936 13874
rect 28172 13388 28224 13394
rect 28172 13330 28224 13336
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27896 13320 27948 13326
rect 27896 13262 27948 13268
rect 27816 12918 27844 13262
rect 27896 13184 27948 13190
rect 27896 13126 27948 13132
rect 27804 12912 27856 12918
rect 27804 12854 27856 12860
rect 27724 12406 27844 12434
rect 27620 11756 27672 11762
rect 27672 11716 27752 11744
rect 27620 11698 27672 11704
rect 27528 11280 27580 11286
rect 27528 11222 27580 11228
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27528 11076 27580 11082
rect 27528 11018 27580 11024
rect 27540 10810 27568 11018
rect 27528 10804 27580 10810
rect 27528 10746 27580 10752
rect 27632 9450 27660 11086
rect 27724 10742 27752 11716
rect 27712 10736 27764 10742
rect 27712 10678 27764 10684
rect 27620 9444 27672 9450
rect 27620 9386 27672 9392
rect 27448 9302 27568 9330
rect 27344 9172 27396 9178
rect 27344 9114 27396 9120
rect 27436 9172 27488 9178
rect 27436 9114 27488 9120
rect 27448 8362 27476 9114
rect 27540 8634 27568 9302
rect 27528 8628 27580 8634
rect 27528 8570 27580 8576
rect 27436 8356 27488 8362
rect 27436 8298 27488 8304
rect 27448 7886 27476 8298
rect 27436 7880 27488 7886
rect 27436 7822 27488 7828
rect 27540 7818 27568 8570
rect 27528 7812 27580 7818
rect 27528 7754 27580 7760
rect 26976 7744 27028 7750
rect 26976 7686 27028 7692
rect 27816 7410 27844 12406
rect 27908 10198 27936 13126
rect 28080 12436 28132 12442
rect 28080 12378 28132 12384
rect 28092 12170 28120 12378
rect 28184 12238 28212 13330
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28080 12164 28132 12170
rect 28080 12106 28132 12112
rect 27988 11892 28040 11898
rect 27988 11834 28040 11840
rect 28000 11014 28028 11834
rect 28092 11150 28120 12106
rect 28080 11144 28132 11150
rect 28080 11086 28132 11092
rect 27988 11008 28040 11014
rect 27988 10950 28040 10956
rect 27896 10192 27948 10198
rect 27896 10134 27948 10140
rect 28000 10062 28028 10950
rect 27988 10056 28040 10062
rect 27988 9998 28040 10004
rect 28172 9920 28224 9926
rect 28172 9862 28224 9868
rect 28184 8974 28212 9862
rect 28264 9716 28316 9722
rect 28264 9658 28316 9664
rect 28276 9042 28304 9658
rect 28264 9036 28316 9042
rect 28264 8978 28316 8984
rect 28172 8968 28224 8974
rect 28172 8910 28224 8916
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 27804 7404 27856 7410
rect 27804 7346 27856 7352
rect 26884 6996 26936 7002
rect 26884 6938 26936 6944
rect 27816 6882 27844 7346
rect 28276 7206 28304 7754
rect 28264 7200 28316 7206
rect 28264 7142 28316 7148
rect 26976 6860 27028 6866
rect 27816 6854 27936 6882
rect 26976 6802 27028 6808
rect 26988 5846 27016 6802
rect 27908 6798 27936 6854
rect 27896 6792 27948 6798
rect 27896 6734 27948 6740
rect 28276 6730 28304 7142
rect 28264 6724 28316 6730
rect 28264 6666 28316 6672
rect 26976 5840 27028 5846
rect 26976 5782 27028 5788
rect 26792 5568 26844 5574
rect 26792 5510 26844 5516
rect 28368 4078 28396 16351
rect 28460 16182 28488 17070
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28460 15502 28488 16118
rect 28448 15496 28500 15502
rect 28448 15438 28500 15444
rect 28552 14498 28580 32846
rect 28632 32428 28684 32434
rect 28632 32370 28684 32376
rect 28644 32230 28672 32370
rect 28632 32224 28684 32230
rect 28632 32166 28684 32172
rect 28632 27328 28684 27334
rect 28630 27296 28632 27305
rect 28684 27296 28686 27305
rect 28630 27231 28686 27240
rect 28736 22094 28764 35006
rect 28828 31414 28856 39238
rect 28908 38344 28960 38350
rect 28908 38286 28960 38292
rect 29012 38298 29040 39374
rect 29092 38344 29144 38350
rect 29012 38292 29092 38298
rect 29012 38286 29144 38292
rect 28920 38214 28948 38286
rect 29012 38270 29132 38286
rect 28908 38208 28960 38214
rect 28908 38150 28960 38156
rect 29012 37942 29040 38270
rect 29000 37936 29052 37942
rect 29000 37878 29052 37884
rect 29184 37868 29236 37874
rect 29184 37810 29236 37816
rect 29000 34672 29052 34678
rect 29000 34614 29052 34620
rect 29012 33946 29040 34614
rect 29196 34406 29224 37810
rect 29184 34400 29236 34406
rect 29184 34342 29236 34348
rect 28920 33918 29040 33946
rect 29092 33924 29144 33930
rect 28920 33522 28948 33918
rect 29092 33866 29144 33872
rect 29000 33856 29052 33862
rect 29000 33798 29052 33804
rect 28908 33516 28960 33522
rect 28908 33458 28960 33464
rect 29012 32994 29040 33798
rect 29104 33046 29132 33866
rect 28920 32966 29040 32994
rect 29092 33040 29144 33046
rect 29092 32982 29144 32988
rect 28920 32910 28948 32966
rect 28908 32904 28960 32910
rect 28908 32846 28960 32852
rect 29000 32904 29052 32910
rect 29000 32846 29052 32852
rect 29012 32434 29040 32846
rect 29184 32836 29236 32842
rect 29184 32778 29236 32784
rect 29000 32428 29052 32434
rect 29000 32370 29052 32376
rect 28908 32292 28960 32298
rect 28908 32234 28960 32240
rect 28920 31890 28948 32234
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28816 31408 28868 31414
rect 28816 31350 28868 31356
rect 28920 31210 28948 31826
rect 29092 31680 29144 31686
rect 29092 31622 29144 31628
rect 28908 31204 28960 31210
rect 28908 31146 28960 31152
rect 29104 30598 29132 31622
rect 29196 31142 29224 32778
rect 29184 31136 29236 31142
rect 29184 31078 29236 31084
rect 29196 30734 29224 31078
rect 29184 30728 29236 30734
rect 29184 30670 29236 30676
rect 29092 30592 29144 30598
rect 29092 30534 29144 30540
rect 29184 30592 29236 30598
rect 29184 30534 29236 30540
rect 29104 30394 29132 30534
rect 29092 30388 29144 30394
rect 29092 30330 29144 30336
rect 29000 29232 29052 29238
rect 29000 29174 29052 29180
rect 29012 28694 29040 29174
rect 29196 29170 29224 30534
rect 29288 30297 29316 48622
rect 29564 48346 29592 48622
rect 29552 48340 29604 48346
rect 29552 48282 29604 48288
rect 29552 48136 29604 48142
rect 29552 48078 29604 48084
rect 29564 47190 29592 48078
rect 29552 47184 29604 47190
rect 29552 47126 29604 47132
rect 29828 40724 29880 40730
rect 29828 40666 29880 40672
rect 29840 39302 29868 40666
rect 29828 39296 29880 39302
rect 29828 39238 29880 39244
rect 29368 37868 29420 37874
rect 29368 37810 29420 37816
rect 29380 36922 29408 37810
rect 29644 37664 29696 37670
rect 29644 37606 29696 37612
rect 29656 37262 29684 37606
rect 29644 37256 29696 37262
rect 29644 37198 29696 37204
rect 29644 37120 29696 37126
rect 29644 37062 29696 37068
rect 29368 36916 29420 36922
rect 29368 36858 29420 36864
rect 29656 36582 29684 37062
rect 29840 36786 29868 39238
rect 29828 36780 29880 36786
rect 29828 36722 29880 36728
rect 29644 36576 29696 36582
rect 29644 36518 29696 36524
rect 29460 34604 29512 34610
rect 29460 34546 29512 34552
rect 29368 33516 29420 33522
rect 29368 33458 29420 33464
rect 29380 33046 29408 33458
rect 29368 33040 29420 33046
rect 29368 32982 29420 32988
rect 29472 32842 29500 34546
rect 29552 33992 29604 33998
rect 29552 33934 29604 33940
rect 29564 33590 29592 33934
rect 29552 33584 29604 33590
rect 29552 33526 29604 33532
rect 29460 32836 29512 32842
rect 29460 32778 29512 32784
rect 29656 32366 29684 36518
rect 29736 34604 29788 34610
rect 29736 34546 29788 34552
rect 29748 32910 29776 34546
rect 29828 33448 29880 33454
rect 29828 33390 29880 33396
rect 29840 32978 29868 33390
rect 29828 32972 29880 32978
rect 29828 32914 29880 32920
rect 29736 32904 29788 32910
rect 29736 32846 29788 32852
rect 29840 32366 29868 32914
rect 29644 32360 29696 32366
rect 29644 32302 29696 32308
rect 29828 32360 29880 32366
rect 29828 32302 29880 32308
rect 29736 32020 29788 32026
rect 29736 31962 29788 31968
rect 29748 31754 29776 31962
rect 29840 31890 29868 32302
rect 29828 31884 29880 31890
rect 29828 31826 29880 31832
rect 29552 31748 29604 31754
rect 29552 31690 29604 31696
rect 29736 31748 29788 31754
rect 29736 31690 29788 31696
rect 29564 31482 29592 31690
rect 29552 31476 29604 31482
rect 29552 31418 29604 31424
rect 29644 31340 29696 31346
rect 29644 31282 29696 31288
rect 29274 30288 29330 30297
rect 29274 30223 29330 30232
rect 29288 30190 29316 30223
rect 29276 30184 29328 30190
rect 29276 30126 29328 30132
rect 29656 29306 29684 31282
rect 29736 31272 29788 31278
rect 29736 31214 29788 31220
rect 29644 29300 29696 29306
rect 29644 29242 29696 29248
rect 29368 29232 29420 29238
rect 29288 29192 29368 29220
rect 29184 29164 29236 29170
rect 29184 29106 29236 29112
rect 29000 28688 29052 28694
rect 29000 28630 29052 28636
rect 29288 28121 29316 29192
rect 29368 29174 29420 29180
rect 29552 28688 29604 28694
rect 29552 28630 29604 28636
rect 29368 28484 29420 28490
rect 29368 28426 29420 28432
rect 29274 28112 29330 28121
rect 29274 28047 29276 28056
rect 29328 28047 29330 28056
rect 29276 28018 29328 28024
rect 28908 28008 28960 28014
rect 28908 27950 28960 27956
rect 28920 27062 28948 27950
rect 29000 27872 29052 27878
rect 29000 27814 29052 27820
rect 29012 27470 29040 27814
rect 29000 27464 29052 27470
rect 29000 27406 29052 27412
rect 29184 27328 29236 27334
rect 29184 27270 29236 27276
rect 29196 27062 29224 27270
rect 28908 27056 28960 27062
rect 28908 26998 28960 27004
rect 29184 27056 29236 27062
rect 29184 26998 29236 27004
rect 29196 25906 29224 26998
rect 29380 26994 29408 28426
rect 29564 27538 29592 28630
rect 29644 28076 29696 28082
rect 29644 28018 29696 28024
rect 29552 27532 29604 27538
rect 29552 27474 29604 27480
rect 29656 27130 29684 28018
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29368 26988 29420 26994
rect 29368 26930 29420 26936
rect 29552 26852 29604 26858
rect 29552 26794 29604 26800
rect 29564 26761 29592 26794
rect 29644 26784 29696 26790
rect 29550 26752 29606 26761
rect 29644 26726 29696 26732
rect 29550 26687 29606 26696
rect 29656 25974 29684 26726
rect 29644 25968 29696 25974
rect 29644 25910 29696 25916
rect 29184 25900 29236 25906
rect 29184 25842 29236 25848
rect 28816 25492 28868 25498
rect 28816 25434 28868 25440
rect 28828 25226 28856 25434
rect 29644 25288 29696 25294
rect 29644 25230 29696 25236
rect 28816 25220 28868 25226
rect 28816 25162 28868 25168
rect 28908 25220 28960 25226
rect 28908 25162 28960 25168
rect 28920 24041 28948 25162
rect 29552 24744 29604 24750
rect 29552 24686 29604 24692
rect 29092 24268 29144 24274
rect 29092 24210 29144 24216
rect 29000 24064 29052 24070
rect 28906 24032 28962 24041
rect 29104 24052 29132 24210
rect 29052 24024 29132 24052
rect 29000 24006 29052 24012
rect 28906 23967 28962 23976
rect 28908 23588 28960 23594
rect 28908 23530 28960 23536
rect 28920 23186 28948 23530
rect 28908 23180 28960 23186
rect 28908 23122 28960 23128
rect 28736 22066 28856 22094
rect 28724 20868 28776 20874
rect 28724 20810 28776 20816
rect 28632 19780 28684 19786
rect 28632 19722 28684 19728
rect 28644 19514 28672 19722
rect 28632 19508 28684 19514
rect 28632 19450 28684 19456
rect 28632 19236 28684 19242
rect 28632 19178 28684 19184
rect 28644 18698 28672 19178
rect 28736 18834 28764 20810
rect 28724 18828 28776 18834
rect 28724 18770 28776 18776
rect 28632 18692 28684 18698
rect 28632 18634 28684 18640
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28736 17270 28764 17478
rect 28724 17264 28776 17270
rect 28724 17206 28776 17212
rect 28724 16516 28776 16522
rect 28724 16458 28776 16464
rect 28736 15502 28764 16458
rect 28724 15496 28776 15502
rect 28724 15438 28776 15444
rect 28552 14470 28764 14498
rect 28632 11620 28684 11626
rect 28632 11562 28684 11568
rect 28644 11150 28672 11562
rect 28632 11144 28684 11150
rect 28632 11086 28684 11092
rect 28448 11008 28500 11014
rect 28448 10950 28500 10956
rect 28460 10130 28488 10950
rect 28540 10192 28592 10198
rect 28540 10134 28592 10140
rect 28448 10124 28500 10130
rect 28448 10066 28500 10072
rect 28552 9518 28580 10134
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28448 9512 28500 9518
rect 28448 9454 28500 9460
rect 28540 9512 28592 9518
rect 28540 9454 28592 9460
rect 28460 9042 28488 9454
rect 28540 9104 28592 9110
rect 28540 9046 28592 9052
rect 28448 9036 28500 9042
rect 28448 8978 28500 8984
rect 28552 8974 28580 9046
rect 28644 8974 28672 9522
rect 28540 8968 28592 8974
rect 28540 8910 28592 8916
rect 28632 8968 28684 8974
rect 28632 8910 28684 8916
rect 28356 4072 28408 4078
rect 28356 4014 28408 4020
rect 26700 3188 26752 3194
rect 26700 3130 26752 3136
rect 26712 2990 26740 3130
rect 26700 2984 26752 2990
rect 26700 2926 26752 2932
rect 27252 2576 27304 2582
rect 27252 2518 27304 2524
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 26516 1896 26568 1902
rect 26516 1838 26568 1844
rect 27080 800 27108 2382
rect 27264 2106 27292 2518
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 27252 2100 27304 2106
rect 27252 2042 27304 2048
rect 27724 800 27752 2382
rect 28736 1970 28764 14470
rect 28828 8906 28856 22066
rect 28920 21554 28948 23122
rect 29012 23118 29040 24006
rect 29368 23724 29420 23730
rect 29368 23666 29420 23672
rect 29092 23180 29144 23186
rect 29092 23122 29144 23128
rect 29000 23112 29052 23118
rect 29000 23054 29052 23060
rect 29104 22166 29132 23122
rect 29380 23050 29408 23666
rect 29564 23526 29592 24686
rect 29656 24206 29684 25230
rect 29748 24614 29776 31214
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 29840 28150 29868 29242
rect 29828 28144 29880 28150
rect 29828 28086 29880 28092
rect 29736 24608 29788 24614
rect 29736 24550 29788 24556
rect 29644 24200 29696 24206
rect 29644 24142 29696 24148
rect 29552 23520 29604 23526
rect 29552 23462 29604 23468
rect 29828 23112 29880 23118
rect 29828 23054 29880 23060
rect 29368 23044 29420 23050
rect 29368 22986 29420 22992
rect 29092 22160 29144 22166
rect 29092 22102 29144 22108
rect 29380 21622 29408 22986
rect 29840 22710 29868 23054
rect 29828 22704 29880 22710
rect 29828 22646 29880 22652
rect 29460 22636 29512 22642
rect 29460 22578 29512 22584
rect 29736 22636 29788 22642
rect 29736 22578 29788 22584
rect 29472 22438 29500 22578
rect 29460 22432 29512 22438
rect 29460 22374 29512 22380
rect 29184 21616 29236 21622
rect 29184 21558 29236 21564
rect 29368 21616 29420 21622
rect 29368 21558 29420 21564
rect 28908 21548 28960 21554
rect 28908 21490 28960 21496
rect 28908 19372 28960 19378
rect 28908 19314 28960 19320
rect 29092 19372 29144 19378
rect 29092 19314 29144 19320
rect 28920 18902 28948 19314
rect 29104 18970 29132 19314
rect 29092 18964 29144 18970
rect 29092 18906 29144 18912
rect 28908 18896 28960 18902
rect 28908 18838 28960 18844
rect 29000 18080 29052 18086
rect 29000 18022 29052 18028
rect 29012 17610 29040 18022
rect 29196 17746 29224 21558
rect 29472 21078 29500 22374
rect 29748 22234 29776 22578
rect 29736 22228 29788 22234
rect 29736 22170 29788 22176
rect 29552 22024 29604 22030
rect 29552 21966 29604 21972
rect 29564 21894 29592 21966
rect 29552 21888 29604 21894
rect 29552 21830 29604 21836
rect 29564 21622 29592 21830
rect 29552 21616 29604 21622
rect 29552 21558 29604 21564
rect 29644 21616 29696 21622
rect 29644 21558 29696 21564
rect 29656 21418 29684 21558
rect 29644 21412 29696 21418
rect 29644 21354 29696 21360
rect 29460 21072 29512 21078
rect 29460 21014 29512 21020
rect 29748 20534 29776 22170
rect 29932 21962 29960 49302
rect 30944 49298 30972 51200
rect 30472 49292 30524 49298
rect 30472 49234 30524 49240
rect 30932 49292 30984 49298
rect 30932 49234 30984 49240
rect 30484 47666 30512 49234
rect 31944 49224 31996 49230
rect 31944 49166 31996 49172
rect 30656 49156 30708 49162
rect 30656 49098 30708 49104
rect 30668 48278 30696 49098
rect 30656 48272 30708 48278
rect 30656 48214 30708 48220
rect 31956 48210 31984 49166
rect 32128 49088 32180 49094
rect 32128 49030 32180 49036
rect 32140 48754 32168 49030
rect 32128 48748 32180 48754
rect 32128 48690 32180 48696
rect 32232 48210 32260 51200
rect 33060 48770 33088 51326
rect 33506 51200 33562 52000
rect 34150 51354 34206 52000
rect 34794 51354 34850 52000
rect 33796 51326 34206 51354
rect 33520 49366 33548 51200
rect 33508 49360 33560 49366
rect 33508 49302 33560 49308
rect 33508 49224 33560 49230
rect 33508 49166 33560 49172
rect 33060 48742 33180 48770
rect 33152 48686 33180 48742
rect 32312 48680 32364 48686
rect 32312 48622 32364 48628
rect 33140 48680 33192 48686
rect 33140 48622 33192 48628
rect 31944 48204 31996 48210
rect 31944 48146 31996 48152
rect 32220 48204 32272 48210
rect 32220 48146 32272 48152
rect 30564 48136 30616 48142
rect 30564 48078 30616 48084
rect 30472 47660 30524 47666
rect 30472 47602 30524 47608
rect 30576 46102 30604 48078
rect 31116 48068 31168 48074
rect 31116 48010 31168 48016
rect 31128 47802 31156 48010
rect 32324 47802 32352 48622
rect 33324 48136 33376 48142
rect 33324 48078 33376 48084
rect 31116 47796 31168 47802
rect 31116 47738 31168 47744
rect 32312 47796 32364 47802
rect 32312 47738 32364 47744
rect 31024 47660 31076 47666
rect 31024 47602 31076 47608
rect 32404 47660 32456 47666
rect 32404 47602 32456 47608
rect 31036 47462 31064 47602
rect 31024 47456 31076 47462
rect 31024 47398 31076 47404
rect 31300 47456 31352 47462
rect 31300 47398 31352 47404
rect 30564 46096 30616 46102
rect 30564 46038 30616 46044
rect 30932 37120 30984 37126
rect 30932 37062 30984 37068
rect 30944 36786 30972 37062
rect 30012 36780 30064 36786
rect 30012 36722 30064 36728
rect 30932 36780 30984 36786
rect 30932 36722 30984 36728
rect 30024 36310 30052 36722
rect 30012 36304 30064 36310
rect 30012 36246 30064 36252
rect 30104 34604 30156 34610
rect 30104 34546 30156 34552
rect 30012 32768 30064 32774
rect 30012 32710 30064 32716
rect 30024 32570 30052 32710
rect 30012 32564 30064 32570
rect 30012 32506 30064 32512
rect 30116 32366 30144 34546
rect 30380 34536 30432 34542
rect 30380 34478 30432 34484
rect 30392 33522 30420 34478
rect 31208 34196 31260 34202
rect 31208 34138 31260 34144
rect 31220 33998 31248 34138
rect 31208 33992 31260 33998
rect 31208 33934 31260 33940
rect 30932 33856 30984 33862
rect 30932 33798 30984 33804
rect 30944 33658 30972 33798
rect 30932 33652 30984 33658
rect 30932 33594 30984 33600
rect 30380 33516 30432 33522
rect 30380 33458 30432 33464
rect 31220 33386 31248 33934
rect 31208 33380 31260 33386
rect 31208 33322 31260 33328
rect 30288 32836 30340 32842
rect 30288 32778 30340 32784
rect 30104 32360 30156 32366
rect 30104 32302 30156 32308
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 30024 30734 30052 31622
rect 30012 30728 30064 30734
rect 30012 30670 30064 30676
rect 30116 28626 30144 32302
rect 30196 32224 30248 32230
rect 30196 32166 30248 32172
rect 30208 31346 30236 32166
rect 30300 31906 30328 32778
rect 30300 31878 30420 31906
rect 30392 31362 30420 31878
rect 30472 31748 30524 31754
rect 30472 31690 30524 31696
rect 30484 31482 30512 31690
rect 30472 31476 30524 31482
rect 30472 31418 30524 31424
rect 30300 31346 30420 31362
rect 30196 31340 30248 31346
rect 30196 31282 30248 31288
rect 30300 31340 30432 31346
rect 30300 31334 30380 31340
rect 30196 31204 30248 31210
rect 30196 31146 30248 31152
rect 30208 30938 30236 31146
rect 30196 30932 30248 30938
rect 30196 30874 30248 30880
rect 30300 30734 30328 31334
rect 30380 31282 30432 31288
rect 30932 31340 30984 31346
rect 30932 31282 30984 31288
rect 30288 30728 30340 30734
rect 30288 30670 30340 30676
rect 30944 30258 30972 31282
rect 30932 30252 30984 30258
rect 30932 30194 30984 30200
rect 30944 29646 30972 30194
rect 31208 29708 31260 29714
rect 31208 29650 31260 29656
rect 30932 29640 30984 29646
rect 30932 29582 30984 29588
rect 30840 28960 30892 28966
rect 30840 28902 30892 28908
rect 30104 28620 30156 28626
rect 30104 28562 30156 28568
rect 30852 28558 30880 28902
rect 31220 28626 31248 29650
rect 31208 28620 31260 28626
rect 31208 28562 31260 28568
rect 30840 28552 30892 28558
rect 30840 28494 30892 28500
rect 30380 28076 30432 28082
rect 30380 28018 30432 28024
rect 30392 26994 30420 28018
rect 31312 28014 31340 47398
rect 32416 47122 32444 47602
rect 32404 47116 32456 47122
rect 32404 47058 32456 47064
rect 33232 47116 33284 47122
rect 33232 47058 33284 47064
rect 31668 46096 31720 46102
rect 31668 46038 31720 46044
rect 31484 33312 31536 33318
rect 31484 33254 31536 33260
rect 31496 32910 31524 33254
rect 31484 32904 31536 32910
rect 31484 32846 31536 32852
rect 31680 30682 31708 46038
rect 33048 37324 33100 37330
rect 33048 37266 33100 37272
rect 32312 35080 32364 35086
rect 32312 35022 32364 35028
rect 32324 34746 32352 35022
rect 32312 34740 32364 34746
rect 32312 34682 32364 34688
rect 31760 34604 31812 34610
rect 31760 34546 31812 34552
rect 31772 34202 31800 34546
rect 31944 34536 31996 34542
rect 31944 34478 31996 34484
rect 32128 34536 32180 34542
rect 32128 34478 32180 34484
rect 31760 34196 31812 34202
rect 31760 34138 31812 34144
rect 31956 33998 31984 34478
rect 31944 33992 31996 33998
rect 31944 33934 31996 33940
rect 32140 33930 32168 34478
rect 32404 34060 32456 34066
rect 32404 34002 32456 34008
rect 32128 33924 32180 33930
rect 32128 33866 32180 33872
rect 31760 33856 31812 33862
rect 31760 33798 31812 33804
rect 31772 33590 31800 33798
rect 31760 33584 31812 33590
rect 31760 33526 31812 33532
rect 31772 32298 31800 33526
rect 32416 33504 32444 34002
rect 32588 33924 32640 33930
rect 32588 33866 32640 33872
rect 32600 33658 32628 33866
rect 32588 33652 32640 33658
rect 32588 33594 32640 33600
rect 32588 33516 32640 33522
rect 32416 33476 32588 33504
rect 32588 33458 32640 33464
rect 32772 33516 32824 33522
rect 32772 33458 32824 33464
rect 32404 32836 32456 32842
rect 32404 32778 32456 32784
rect 32416 32434 32444 32778
rect 31852 32428 31904 32434
rect 31852 32370 31904 32376
rect 32404 32428 32456 32434
rect 32404 32370 32456 32376
rect 31760 32292 31812 32298
rect 31760 32234 31812 32240
rect 31772 31822 31800 32234
rect 31864 32026 31892 32370
rect 31852 32020 31904 32026
rect 31852 31962 31904 31968
rect 31760 31816 31812 31822
rect 31760 31758 31812 31764
rect 31496 30654 31708 30682
rect 31392 30388 31444 30394
rect 31392 30330 31444 30336
rect 31404 29578 31432 30330
rect 31392 29572 31444 29578
rect 31392 29514 31444 29520
rect 31404 29170 31432 29514
rect 31392 29164 31444 29170
rect 31392 29106 31444 29112
rect 31496 29050 31524 30654
rect 31668 30592 31720 30598
rect 31668 30534 31720 30540
rect 31680 30258 31708 30534
rect 31668 30252 31720 30258
rect 31668 30194 31720 30200
rect 31680 29782 31708 30194
rect 31668 29776 31720 29782
rect 31668 29718 31720 29724
rect 31772 29714 31800 31758
rect 31864 31414 31892 31962
rect 32128 31748 32180 31754
rect 32128 31690 32180 31696
rect 32140 31482 32168 31690
rect 32128 31476 32180 31482
rect 32128 31418 32180 31424
rect 31852 31408 31904 31414
rect 31852 31350 31904 31356
rect 32600 31346 32628 33458
rect 32784 33114 32812 33458
rect 32772 33108 32824 33114
rect 32772 33050 32824 33056
rect 32772 32224 32824 32230
rect 32772 32166 32824 32172
rect 32784 31346 32812 32166
rect 33060 31754 33088 37266
rect 32876 31726 33088 31754
rect 32588 31340 32640 31346
rect 32508 31300 32588 31328
rect 32220 30592 32272 30598
rect 32220 30534 32272 30540
rect 31944 30252 31996 30258
rect 31944 30194 31996 30200
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31956 30054 31984 30194
rect 31852 30048 31904 30054
rect 31852 29990 31904 29996
rect 31944 30048 31996 30054
rect 31944 29990 31996 29996
rect 31760 29708 31812 29714
rect 31760 29650 31812 29656
rect 31772 29170 31800 29650
rect 31864 29646 31892 29990
rect 32140 29850 32168 30194
rect 32128 29844 32180 29850
rect 32128 29786 32180 29792
rect 31852 29640 31904 29646
rect 31852 29582 31904 29588
rect 32232 29578 32260 30534
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32324 30054 32352 30194
rect 32312 30048 32364 30054
rect 32312 29990 32364 29996
rect 32220 29572 32272 29578
rect 32220 29514 32272 29520
rect 32128 29504 32180 29510
rect 32128 29446 32180 29452
rect 32140 29238 32168 29446
rect 32128 29232 32180 29238
rect 32324 29186 32352 29990
rect 32128 29174 32180 29180
rect 31760 29164 31812 29170
rect 31760 29106 31812 29112
rect 32232 29158 32352 29186
rect 31404 29022 31524 29050
rect 32128 29096 32180 29102
rect 32128 29038 32180 29044
rect 30748 28008 30800 28014
rect 30748 27950 30800 27956
rect 31300 28008 31352 28014
rect 31300 27950 31352 27956
rect 30564 27532 30616 27538
rect 30564 27474 30616 27480
rect 30576 27062 30604 27474
rect 30564 27056 30616 27062
rect 30564 26998 30616 27004
rect 30380 26988 30432 26994
rect 30380 26930 30432 26936
rect 30392 26314 30420 26930
rect 30472 26920 30524 26926
rect 30472 26862 30524 26868
rect 30380 26308 30432 26314
rect 30380 26250 30432 26256
rect 30484 26246 30512 26862
rect 30472 26240 30524 26246
rect 30472 26182 30524 26188
rect 30012 24132 30064 24138
rect 30012 24074 30064 24080
rect 30024 23866 30052 24074
rect 30012 23860 30064 23866
rect 30012 23802 30064 23808
rect 30380 23860 30432 23866
rect 30380 23802 30432 23808
rect 30024 22094 30052 23802
rect 30392 23746 30420 23802
rect 30300 23730 30420 23746
rect 30288 23724 30420 23730
rect 30340 23718 30420 23724
rect 30472 23724 30524 23730
rect 30288 23666 30340 23672
rect 30472 23666 30524 23672
rect 30196 23656 30248 23662
rect 30196 23598 30248 23604
rect 30208 22642 30236 23598
rect 30380 23520 30432 23526
rect 30380 23462 30432 23468
rect 30392 23118 30420 23462
rect 30484 23322 30512 23666
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30656 23112 30708 23118
rect 30656 23054 30708 23060
rect 30564 22772 30616 22778
rect 30564 22714 30616 22720
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30024 22066 30144 22094
rect 29920 21956 29972 21962
rect 29920 21898 29972 21904
rect 29276 20528 29328 20534
rect 29276 20470 29328 20476
rect 29736 20528 29788 20534
rect 29736 20470 29788 20476
rect 29288 19378 29316 20470
rect 30012 19712 30064 19718
rect 30012 19654 30064 19660
rect 30024 19378 30052 19654
rect 29276 19372 29328 19378
rect 30012 19372 30064 19378
rect 29276 19314 29328 19320
rect 29932 19320 30012 19334
rect 29932 19314 30064 19320
rect 29932 19306 30052 19314
rect 29932 18698 29960 19306
rect 29920 18692 29972 18698
rect 29920 18634 29972 18640
rect 29276 18624 29328 18630
rect 29276 18566 29328 18572
rect 29184 17740 29236 17746
rect 29184 17682 29236 17688
rect 29288 17678 29316 18566
rect 29276 17672 29328 17678
rect 29276 17614 29328 17620
rect 29000 17604 29052 17610
rect 29000 17546 29052 17552
rect 28908 17196 28960 17202
rect 28908 17138 28960 17144
rect 28920 15706 28948 17138
rect 29012 16674 29040 17546
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29196 16998 29224 17138
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29012 16658 29132 16674
rect 29012 16652 29144 16658
rect 29012 16646 29092 16652
rect 29092 16594 29144 16600
rect 29000 16244 29052 16250
rect 29000 16186 29052 16192
rect 28908 15700 28960 15706
rect 28908 15642 28960 15648
rect 29012 15094 29040 16186
rect 29196 16182 29224 16934
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29184 15904 29236 15910
rect 29184 15846 29236 15852
rect 29000 15088 29052 15094
rect 29000 15030 29052 15036
rect 29196 14074 29224 15846
rect 29288 14414 29316 17614
rect 29828 17536 29880 17542
rect 29828 17478 29880 17484
rect 29460 17264 29512 17270
rect 29460 17206 29512 17212
rect 29472 16114 29500 17206
rect 29736 16992 29788 16998
rect 29736 16934 29788 16940
rect 29748 16726 29776 16934
rect 29736 16720 29788 16726
rect 29736 16662 29788 16668
rect 29840 16590 29868 17478
rect 29828 16584 29880 16590
rect 29828 16526 29880 16532
rect 29736 16516 29788 16522
rect 29736 16458 29788 16464
rect 29460 16108 29512 16114
rect 29460 16050 29512 16056
rect 29472 15366 29500 16050
rect 29552 16040 29604 16046
rect 29552 15982 29604 15988
rect 29564 15881 29592 15982
rect 29550 15872 29606 15881
rect 29550 15807 29606 15816
rect 29644 15428 29696 15434
rect 29644 15370 29696 15376
rect 29460 15360 29512 15366
rect 29460 15302 29512 15308
rect 29656 15026 29684 15370
rect 29644 15020 29696 15026
rect 29644 14962 29696 14968
rect 29552 14952 29604 14958
rect 29552 14894 29604 14900
rect 29368 14816 29420 14822
rect 29368 14758 29420 14764
rect 29460 14816 29512 14822
rect 29460 14758 29512 14764
rect 29380 14550 29408 14758
rect 29368 14544 29420 14550
rect 29368 14486 29420 14492
rect 29276 14408 29328 14414
rect 29276 14350 29328 14356
rect 29184 14068 29236 14074
rect 29184 14010 29236 14016
rect 29288 13326 29316 14350
rect 29380 13530 29408 14486
rect 29472 13938 29500 14758
rect 29564 14618 29592 14894
rect 29552 14612 29604 14618
rect 29552 14554 29604 14560
rect 29656 13938 29684 14962
rect 29460 13932 29512 13938
rect 29460 13874 29512 13880
rect 29644 13932 29696 13938
rect 29644 13874 29696 13880
rect 29368 13524 29420 13530
rect 29368 13466 29420 13472
rect 29472 13462 29500 13874
rect 29656 13818 29684 13874
rect 29564 13790 29684 13818
rect 29460 13456 29512 13462
rect 29460 13398 29512 13404
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29472 11898 29500 13398
rect 29564 12170 29592 13790
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29656 12850 29684 13126
rect 29644 12844 29696 12850
rect 29644 12786 29696 12792
rect 29748 12782 29776 16458
rect 29828 12844 29880 12850
rect 29828 12786 29880 12792
rect 29736 12776 29788 12782
rect 29736 12718 29788 12724
rect 29840 12442 29868 12786
rect 29828 12436 29880 12442
rect 29828 12378 29880 12384
rect 29644 12300 29696 12306
rect 29644 12242 29696 12248
rect 29552 12164 29604 12170
rect 29552 12106 29604 12112
rect 29460 11892 29512 11898
rect 29460 11834 29512 11840
rect 29276 11756 29328 11762
rect 29276 11698 29328 11704
rect 28908 11552 28960 11558
rect 28960 11512 29040 11540
rect 28908 11494 28960 11500
rect 29012 11121 29040 11512
rect 29288 11354 29316 11698
rect 29656 11694 29684 12242
rect 29828 12232 29880 12238
rect 29828 12174 29880 12180
rect 29644 11688 29696 11694
rect 29644 11630 29696 11636
rect 29552 11620 29604 11626
rect 29552 11562 29604 11568
rect 29276 11348 29328 11354
rect 29276 11290 29328 11296
rect 28998 11112 29054 11121
rect 28998 11047 29054 11056
rect 29564 11014 29592 11562
rect 29552 11008 29604 11014
rect 29552 10950 29604 10956
rect 29368 10804 29420 10810
rect 29012 10764 29368 10792
rect 28908 10736 28960 10742
rect 29012 10724 29040 10764
rect 29368 10746 29420 10752
rect 28960 10696 29040 10724
rect 29460 10736 29512 10742
rect 28908 10678 28960 10684
rect 29460 10678 29512 10684
rect 29276 10668 29328 10674
rect 29276 10610 29328 10616
rect 28998 10432 29054 10441
rect 28998 10367 29054 10376
rect 28908 10056 28960 10062
rect 28906 10024 28908 10033
rect 28960 10024 28962 10033
rect 28906 9959 28962 9968
rect 29012 9586 29040 10367
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 29288 9042 29316 10610
rect 29368 10464 29420 10470
rect 29366 10432 29368 10441
rect 29420 10432 29422 10441
rect 29366 10367 29422 10376
rect 29472 9722 29500 10678
rect 29564 10062 29592 10950
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29552 10056 29604 10062
rect 29552 9998 29604 10004
rect 29748 9722 29776 10610
rect 29840 10266 29868 12174
rect 29932 11150 29960 18634
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30024 17338 30052 17682
rect 30116 17490 30144 22066
rect 30208 20466 30236 22578
rect 30576 21690 30604 22714
rect 30668 22166 30696 23054
rect 30656 22160 30708 22166
rect 30656 22102 30708 22108
rect 30564 21684 30616 21690
rect 30564 21626 30616 21632
rect 30656 20868 30708 20874
rect 30656 20810 30708 20816
rect 30196 20460 30248 20466
rect 30196 20402 30248 20408
rect 30288 20460 30340 20466
rect 30288 20402 30340 20408
rect 30208 18970 30236 20402
rect 30300 19514 30328 20402
rect 30668 19514 30696 20810
rect 30760 19854 30788 27950
rect 30840 26580 30892 26586
rect 30840 26522 30892 26528
rect 30852 26450 30880 26522
rect 30840 26444 30892 26450
rect 30840 26386 30892 26392
rect 31024 25832 31076 25838
rect 31024 25774 31076 25780
rect 30932 25492 30984 25498
rect 30932 25434 30984 25440
rect 30944 25158 30972 25434
rect 30932 25152 30984 25158
rect 30932 25094 30984 25100
rect 30944 22982 30972 25094
rect 30932 22976 30984 22982
rect 30932 22918 30984 22924
rect 30840 22772 30892 22778
rect 30840 22714 30892 22720
rect 30852 21554 30880 22714
rect 30840 21548 30892 21554
rect 30840 21490 30892 21496
rect 30748 19848 30800 19854
rect 30748 19790 30800 19796
rect 30288 19508 30340 19514
rect 30288 19450 30340 19456
rect 30656 19508 30708 19514
rect 30656 19450 30708 19456
rect 30196 18964 30248 18970
rect 30196 18906 30248 18912
rect 30116 17462 30236 17490
rect 30012 17332 30064 17338
rect 30012 17274 30064 17280
rect 30104 17128 30156 17134
rect 30104 17070 30156 17076
rect 30012 17060 30064 17066
rect 30012 17002 30064 17008
rect 30024 16590 30052 17002
rect 30012 16584 30064 16590
rect 30012 16526 30064 16532
rect 30116 16522 30144 17070
rect 30104 16516 30156 16522
rect 30104 16458 30156 16464
rect 30208 16402 30236 17462
rect 30288 17128 30340 17134
rect 30288 17070 30340 17076
rect 30116 16374 30236 16402
rect 30010 16008 30066 16017
rect 30010 15943 30066 15952
rect 30024 15638 30052 15943
rect 30012 15632 30064 15638
rect 30012 15574 30064 15580
rect 30012 15496 30064 15502
rect 30012 15438 30064 15444
rect 30024 13802 30052 15438
rect 30116 14498 30144 16374
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30208 15502 30236 16186
rect 30300 16017 30328 17070
rect 30564 16244 30616 16250
rect 30564 16186 30616 16192
rect 30286 16008 30342 16017
rect 30286 15943 30342 15952
rect 30380 15904 30432 15910
rect 30380 15846 30432 15852
rect 30288 15700 30340 15706
rect 30288 15642 30340 15648
rect 30196 15496 30248 15502
rect 30196 15438 30248 15444
rect 30300 14890 30328 15642
rect 30392 15162 30420 15846
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30380 15156 30432 15162
rect 30380 15098 30432 15104
rect 30484 15026 30512 15302
rect 30576 15026 30604 16186
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30564 15020 30616 15026
rect 30564 14962 30616 14968
rect 30668 14906 30696 19450
rect 30748 16720 30800 16726
rect 30748 16662 30800 16668
rect 30760 16522 30788 16662
rect 30748 16516 30800 16522
rect 30748 16458 30800 16464
rect 30852 16182 30880 21490
rect 31036 17270 31064 25774
rect 31404 24750 31432 29022
rect 32140 27130 32168 29038
rect 32128 27124 32180 27130
rect 32128 27066 32180 27072
rect 32232 26994 32260 29158
rect 32508 28082 32536 31300
rect 32588 31282 32640 31288
rect 32772 31340 32824 31346
rect 32772 31282 32824 31288
rect 32772 28552 32824 28558
rect 32772 28494 32824 28500
rect 32588 28416 32640 28422
rect 32588 28358 32640 28364
rect 32496 28076 32548 28082
rect 32496 28018 32548 28024
rect 32600 27062 32628 28358
rect 32784 28082 32812 28494
rect 32772 28076 32824 28082
rect 32772 28018 32824 28024
rect 32784 27470 32812 28018
rect 32772 27464 32824 27470
rect 32772 27406 32824 27412
rect 32588 27056 32640 27062
rect 32588 26998 32640 27004
rect 32220 26988 32272 26994
rect 32220 26930 32272 26936
rect 31484 26920 31536 26926
rect 31484 26862 31536 26868
rect 32496 26920 32548 26926
rect 32496 26862 32548 26868
rect 31392 24744 31444 24750
rect 31392 24686 31444 24692
rect 31392 24200 31444 24206
rect 31392 24142 31444 24148
rect 31116 22976 31168 22982
rect 31116 22918 31168 22924
rect 31128 22098 31156 22918
rect 31116 22092 31168 22098
rect 31116 22034 31168 22040
rect 31300 21956 31352 21962
rect 31300 21898 31352 21904
rect 31116 21072 31168 21078
rect 31116 21014 31168 21020
rect 31024 17264 31076 17270
rect 31024 17206 31076 17212
rect 30932 16448 30984 16454
rect 30932 16390 30984 16396
rect 30840 16176 30892 16182
rect 30840 16118 30892 16124
rect 30746 15736 30802 15745
rect 30746 15671 30802 15680
rect 30760 15570 30788 15671
rect 30944 15638 30972 16390
rect 31024 16040 31076 16046
rect 31022 16008 31024 16017
rect 31076 16008 31078 16017
rect 31022 15943 31078 15952
rect 30932 15632 30984 15638
rect 30932 15574 30984 15580
rect 30748 15564 30800 15570
rect 30748 15506 30800 15512
rect 30840 15496 30892 15502
rect 30840 15438 30892 15444
rect 30288 14884 30340 14890
rect 30288 14826 30340 14832
rect 30576 14878 30696 14906
rect 30116 14470 30236 14498
rect 30104 14272 30156 14278
rect 30104 14214 30156 14220
rect 30012 13796 30064 13802
rect 30012 13738 30064 13744
rect 30024 12238 30052 13738
rect 30116 12434 30144 14214
rect 30208 12850 30236 14470
rect 30576 14414 30604 14878
rect 30852 14618 30880 15438
rect 31024 15020 31076 15026
rect 31024 14962 31076 14968
rect 30840 14612 30892 14618
rect 30840 14554 30892 14560
rect 31036 14550 31064 14962
rect 31024 14544 31076 14550
rect 31024 14486 31076 14492
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30840 14408 30892 14414
rect 30840 14350 30892 14356
rect 30656 14340 30708 14346
rect 30656 14282 30708 14288
rect 30668 13870 30696 14282
rect 30656 13864 30708 13870
rect 30656 13806 30708 13812
rect 30668 13326 30696 13806
rect 30748 13796 30800 13802
rect 30748 13738 30800 13744
rect 30656 13320 30708 13326
rect 30656 13262 30708 13268
rect 30564 13184 30616 13190
rect 30564 13126 30616 13132
rect 30196 12844 30248 12850
rect 30196 12786 30248 12792
rect 30576 12434 30604 13126
rect 30656 12912 30708 12918
rect 30656 12854 30708 12860
rect 30116 12406 30236 12434
rect 30012 12232 30064 12238
rect 30012 12174 30064 12180
rect 30104 11620 30156 11626
rect 30104 11562 30156 11568
rect 30116 11218 30144 11562
rect 30104 11212 30156 11218
rect 30104 11154 30156 11160
rect 29920 11144 29972 11150
rect 30208 11098 30236 12406
rect 30484 12406 30604 12434
rect 30484 11762 30512 12406
rect 30472 11756 30524 11762
rect 30472 11698 30524 11704
rect 29920 11086 29972 11092
rect 30116 11070 30236 11098
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 30024 10606 30052 10950
rect 30116 10606 30144 11070
rect 30300 10674 30328 11086
rect 30288 10668 30340 10674
rect 30288 10610 30340 10616
rect 30012 10600 30064 10606
rect 30012 10542 30064 10548
rect 30104 10600 30156 10606
rect 30104 10542 30156 10548
rect 30024 10266 30052 10542
rect 29828 10260 29880 10266
rect 29828 10202 29880 10208
rect 30012 10260 30064 10266
rect 30012 10202 30064 10208
rect 29460 9716 29512 9722
rect 29460 9658 29512 9664
rect 29736 9716 29788 9722
rect 29736 9658 29788 9664
rect 29840 9586 29868 10202
rect 29828 9580 29880 9586
rect 29828 9522 29880 9528
rect 30116 9110 30144 10542
rect 30104 9104 30156 9110
rect 30104 9046 30156 9052
rect 29276 9036 29328 9042
rect 29276 8978 29328 8984
rect 29736 9036 29788 9042
rect 29736 8978 29788 8984
rect 28816 8900 28868 8906
rect 28816 8842 28868 8848
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 28920 8498 28948 8774
rect 29748 8634 29776 8978
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 30484 8498 30512 11698
rect 30668 11694 30696 12854
rect 30760 12714 30788 13738
rect 30852 13734 30880 14350
rect 30932 14068 30984 14074
rect 30932 14010 30984 14016
rect 30944 13870 30972 14010
rect 31024 13932 31076 13938
rect 31024 13874 31076 13880
rect 30932 13864 30984 13870
rect 30932 13806 30984 13812
rect 30840 13728 30892 13734
rect 30840 13670 30892 13676
rect 30748 12708 30800 12714
rect 30748 12650 30800 12656
rect 30760 12170 30788 12650
rect 30840 12640 30892 12646
rect 30840 12582 30892 12588
rect 30748 12164 30800 12170
rect 30748 12106 30800 12112
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 11354 30696 11630
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30564 10668 30616 10674
rect 30564 10610 30616 10616
rect 30576 10198 30604 10610
rect 30668 10538 30696 11290
rect 30760 11218 30788 12106
rect 30748 11212 30800 11218
rect 30748 11154 30800 11160
rect 30656 10532 30708 10538
rect 30656 10474 30708 10480
rect 30564 10192 30616 10198
rect 30760 10146 30788 11154
rect 30852 11150 30880 12582
rect 30840 11144 30892 11150
rect 30840 11086 30892 11092
rect 30944 10674 30972 13806
rect 31036 13530 31064 13874
rect 31024 13524 31076 13530
rect 31024 13466 31076 13472
rect 31128 13190 31156 21014
rect 31208 20936 31260 20942
rect 31208 20878 31260 20884
rect 31220 19990 31248 20878
rect 31208 19984 31260 19990
rect 31208 19926 31260 19932
rect 31116 13184 31168 13190
rect 31116 13126 31168 13132
rect 31312 12434 31340 21898
rect 31404 20330 31432 24142
rect 31392 20324 31444 20330
rect 31392 20266 31444 20272
rect 31404 19922 31432 20266
rect 31392 19916 31444 19922
rect 31392 19858 31444 19864
rect 31392 16516 31444 16522
rect 31392 16458 31444 16464
rect 31404 16114 31432 16458
rect 31392 16108 31444 16114
rect 31392 16050 31444 16056
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31404 14074 31432 14350
rect 31392 14068 31444 14074
rect 31392 14010 31444 14016
rect 31496 12434 31524 26862
rect 32402 26752 32458 26761
rect 32402 26687 32458 26696
rect 32416 26450 32444 26687
rect 32404 26444 32456 26450
rect 32404 26386 32456 26392
rect 31944 26376 31996 26382
rect 31944 26318 31996 26324
rect 31576 25832 31628 25838
rect 31576 25774 31628 25780
rect 31588 23866 31616 25774
rect 31956 25702 31984 26318
rect 32036 25968 32088 25974
rect 32036 25910 32088 25916
rect 31944 25696 31996 25702
rect 31944 25638 31996 25644
rect 31956 24818 31984 25638
rect 32048 24886 32076 25910
rect 32036 24880 32088 24886
rect 32036 24822 32088 24828
rect 31944 24812 31996 24818
rect 31944 24754 31996 24760
rect 31576 23860 31628 23866
rect 31576 23802 31628 23808
rect 32036 22160 32088 22166
rect 32036 22102 32088 22108
rect 31852 21344 31904 21350
rect 31852 21286 31904 21292
rect 31668 20528 31720 20534
rect 31668 20470 31720 20476
rect 31680 19378 31708 20470
rect 31760 19712 31812 19718
rect 31760 19654 31812 19660
rect 31772 19446 31800 19654
rect 31760 19440 31812 19446
rect 31760 19382 31812 19388
rect 31668 19372 31720 19378
rect 31668 19314 31720 19320
rect 31680 17202 31708 19314
rect 31864 18766 31892 21286
rect 32048 20942 32076 22102
rect 32036 20936 32088 20942
rect 32036 20878 32088 20884
rect 32312 20868 32364 20874
rect 32312 20810 32364 20816
rect 32128 20800 32180 20806
rect 32180 20748 32260 20754
rect 32128 20742 32260 20748
rect 32140 20726 32260 20742
rect 32232 20466 32260 20726
rect 32220 20460 32272 20466
rect 32220 20402 32272 20408
rect 32324 19854 32352 20810
rect 32312 19848 32364 19854
rect 32312 19790 32364 19796
rect 32036 19712 32088 19718
rect 32036 19654 32088 19660
rect 31944 19508 31996 19514
rect 31944 19450 31996 19456
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 31864 17898 31892 18702
rect 31956 18630 31984 19450
rect 32048 18766 32076 19654
rect 32416 19514 32444 26386
rect 32508 25906 32536 26862
rect 32496 25900 32548 25906
rect 32496 25842 32548 25848
rect 32496 25696 32548 25702
rect 32496 25638 32548 25644
rect 32508 25294 32536 25638
rect 32496 25288 32548 25294
rect 32496 25230 32548 25236
rect 32496 24812 32548 24818
rect 32496 24754 32548 24760
rect 32508 24342 32536 24754
rect 32588 24744 32640 24750
rect 32588 24686 32640 24692
rect 32496 24336 32548 24342
rect 32496 24278 32548 24284
rect 32508 23730 32536 24278
rect 32496 23724 32548 23730
rect 32496 23666 32548 23672
rect 32508 23118 32536 23666
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32600 20942 32628 24686
rect 32876 24206 32904 31726
rect 33244 30734 33272 47058
rect 33336 35894 33364 48078
rect 33520 47666 33548 49166
rect 33692 48000 33744 48006
rect 33692 47942 33744 47948
rect 33704 47734 33732 47942
rect 33692 47728 33744 47734
rect 33692 47670 33744 47676
rect 33508 47660 33560 47666
rect 33508 47602 33560 47608
rect 33336 35866 33640 35894
rect 33416 35012 33468 35018
rect 33416 34954 33468 34960
rect 33324 33992 33376 33998
rect 33324 33934 33376 33940
rect 33336 33522 33364 33934
rect 33428 33658 33456 34954
rect 33508 34400 33560 34406
rect 33508 34342 33560 34348
rect 33520 33658 33548 34342
rect 33416 33652 33468 33658
rect 33416 33594 33468 33600
rect 33508 33652 33560 33658
rect 33508 33594 33560 33600
rect 33324 33516 33376 33522
rect 33324 33458 33376 33464
rect 33612 31754 33640 35866
rect 33336 31726 33640 31754
rect 33232 30728 33284 30734
rect 33232 30670 33284 30676
rect 33230 30288 33286 30297
rect 33230 30223 33232 30232
rect 33284 30223 33286 30232
rect 33232 30194 33284 30200
rect 33232 28756 33284 28762
rect 33232 28698 33284 28704
rect 33244 28014 33272 28698
rect 33232 28008 33284 28014
rect 33232 27950 33284 27956
rect 33244 26330 33272 27950
rect 33336 26858 33364 31726
rect 33508 30728 33560 30734
rect 33508 30670 33560 30676
rect 33416 30660 33468 30666
rect 33416 30602 33468 30608
rect 33428 29306 33456 30602
rect 33520 29646 33548 30670
rect 33600 30592 33652 30598
rect 33600 30534 33652 30540
rect 33612 30326 33640 30534
rect 33600 30320 33652 30326
rect 33600 30262 33652 30268
rect 33508 29640 33560 29646
rect 33508 29582 33560 29588
rect 33416 29300 33468 29306
rect 33416 29242 33468 29248
rect 33428 28082 33456 29242
rect 33416 28076 33468 28082
rect 33416 28018 33468 28024
rect 33520 27402 33548 29582
rect 33692 29504 33744 29510
rect 33692 29446 33744 29452
rect 33508 27396 33560 27402
rect 33508 27338 33560 27344
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33324 26852 33376 26858
rect 33324 26794 33376 26800
rect 33612 26450 33640 27270
rect 33704 27062 33732 29446
rect 33692 27056 33744 27062
rect 33692 26998 33744 27004
rect 33600 26444 33652 26450
rect 33600 26386 33652 26392
rect 33244 26302 33364 26330
rect 33048 25832 33100 25838
rect 33048 25774 33100 25780
rect 33060 24886 33088 25774
rect 33048 24880 33100 24886
rect 33048 24822 33100 24828
rect 32956 24744 33008 24750
rect 32956 24686 33008 24692
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32968 23866 32996 24686
rect 32956 23860 33008 23866
rect 32956 23802 33008 23808
rect 33232 23656 33284 23662
rect 33232 23598 33284 23604
rect 32680 21956 32732 21962
rect 32680 21898 32732 21904
rect 32864 21956 32916 21962
rect 32864 21898 32916 21904
rect 32692 21486 32720 21898
rect 32680 21480 32732 21486
rect 32680 21422 32732 21428
rect 32692 20942 32720 21422
rect 32876 21350 32904 21898
rect 32864 21344 32916 21350
rect 32864 21286 32916 21292
rect 32588 20936 32640 20942
rect 32588 20878 32640 20884
rect 32680 20936 32732 20942
rect 32680 20878 32732 20884
rect 32600 20482 32628 20878
rect 32600 20466 32720 20482
rect 32600 20460 32732 20466
rect 32600 20454 32680 20460
rect 32680 20402 32732 20408
rect 33244 19854 33272 23598
rect 33336 22094 33364 26302
rect 33508 25356 33560 25362
rect 33508 25298 33560 25304
rect 33520 25158 33548 25298
rect 33692 25288 33744 25294
rect 33692 25230 33744 25236
rect 33704 25158 33732 25230
rect 33508 25152 33560 25158
rect 33508 25094 33560 25100
rect 33692 25152 33744 25158
rect 33692 25094 33744 25100
rect 33704 24342 33732 25094
rect 33692 24336 33744 24342
rect 33692 24278 33744 24284
rect 33704 24206 33732 24278
rect 33692 24200 33744 24206
rect 33692 24142 33744 24148
rect 33416 24064 33468 24070
rect 33416 24006 33468 24012
rect 33428 23662 33456 24006
rect 33796 23662 33824 51326
rect 34150 51200 34206 51326
rect 34716 51326 34850 51354
rect 34428 49360 34480 49366
rect 34428 49302 34480 49308
rect 33876 34536 33928 34542
rect 33876 34478 33928 34484
rect 33888 33862 33916 34478
rect 33968 33992 34020 33998
rect 33968 33934 34020 33940
rect 33876 33856 33928 33862
rect 33876 33798 33928 33804
rect 33888 32910 33916 33798
rect 33876 32904 33928 32910
rect 33876 32846 33928 32852
rect 33876 32496 33928 32502
rect 33876 32438 33928 32444
rect 33888 32026 33916 32438
rect 33876 32020 33928 32026
rect 33876 31962 33928 31968
rect 33980 30734 34008 33934
rect 34336 32020 34388 32026
rect 34336 31962 34388 31968
rect 34348 30734 34376 31962
rect 33968 30728 34020 30734
rect 33968 30670 34020 30676
rect 34336 30728 34388 30734
rect 34336 30670 34388 30676
rect 33980 29646 34008 30670
rect 33968 29640 34020 29646
rect 33968 29582 34020 29588
rect 34060 28960 34112 28966
rect 34060 28902 34112 28908
rect 34072 28490 34100 28902
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 33968 26308 34020 26314
rect 33968 26250 34020 26256
rect 33980 25770 34008 26250
rect 33968 25764 34020 25770
rect 33968 25706 34020 25712
rect 33416 23656 33468 23662
rect 33416 23598 33468 23604
rect 33784 23656 33836 23662
rect 33784 23598 33836 23604
rect 33876 22432 33928 22438
rect 33876 22374 33928 22380
rect 33336 22066 33548 22094
rect 33232 19848 33284 19854
rect 33232 19790 33284 19796
rect 33244 19514 33272 19790
rect 32404 19508 32456 19514
rect 32404 19450 32456 19456
rect 33232 19508 33284 19514
rect 33232 19450 33284 19456
rect 32312 19372 32364 19378
rect 32312 19314 32364 19320
rect 32220 19236 32272 19242
rect 32220 19178 32272 19184
rect 32232 18766 32260 19178
rect 32324 18970 32352 19314
rect 32312 18964 32364 18970
rect 32312 18906 32364 18912
rect 32416 18850 32444 19450
rect 32416 18822 32720 18850
rect 32036 18760 32088 18766
rect 32036 18702 32088 18708
rect 32220 18760 32272 18766
rect 32220 18702 32272 18708
rect 32588 18760 32640 18766
rect 32588 18702 32640 18708
rect 31944 18624 31996 18630
rect 31944 18566 31996 18572
rect 31864 17870 32260 17898
rect 31668 17196 31720 17202
rect 31668 17138 31720 17144
rect 31680 16794 31708 17138
rect 32128 16992 32180 16998
rect 32128 16934 32180 16940
rect 31668 16788 31720 16794
rect 31668 16730 31720 16736
rect 32140 16726 32168 16934
rect 32128 16720 32180 16726
rect 32128 16662 32180 16668
rect 31576 16584 31628 16590
rect 31576 16526 31628 16532
rect 31588 15910 31616 16526
rect 32140 15994 32168 16662
rect 32048 15966 32168 15994
rect 31576 15904 31628 15910
rect 31576 15846 31628 15852
rect 31852 15632 31904 15638
rect 31852 15574 31904 15580
rect 31760 15496 31812 15502
rect 31760 15438 31812 15444
rect 31772 15162 31800 15438
rect 31760 15156 31812 15162
rect 31760 15098 31812 15104
rect 31864 14414 31892 15574
rect 31944 15496 31996 15502
rect 31944 15438 31996 15444
rect 31956 14618 31984 15438
rect 31944 14612 31996 14618
rect 31944 14554 31996 14560
rect 32048 14414 32076 15966
rect 32128 15904 32180 15910
rect 32128 15846 32180 15852
rect 32140 14482 32168 15846
rect 32128 14476 32180 14482
rect 32128 14418 32180 14424
rect 31852 14408 31904 14414
rect 31852 14350 31904 14356
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 32140 14074 32168 14418
rect 32232 14414 32260 17870
rect 32312 16448 32364 16454
rect 32312 16390 32364 16396
rect 32324 16114 32352 16390
rect 32312 16108 32364 16114
rect 32312 16050 32364 16056
rect 32404 16108 32456 16114
rect 32404 16050 32456 16056
rect 32312 15904 32364 15910
rect 32310 15872 32312 15881
rect 32364 15872 32366 15881
rect 32310 15807 32366 15816
rect 32416 15502 32444 16050
rect 32404 15496 32456 15502
rect 32404 15438 32456 15444
rect 32496 15360 32548 15366
rect 32496 15302 32548 15308
rect 32508 15094 32536 15302
rect 32496 15088 32548 15094
rect 32496 15030 32548 15036
rect 32404 14952 32456 14958
rect 32404 14894 32456 14900
rect 32220 14408 32272 14414
rect 32220 14350 32272 14356
rect 32312 14408 32364 14414
rect 32312 14350 32364 14356
rect 32128 14068 32180 14074
rect 32128 14010 32180 14016
rect 32140 13394 32168 14010
rect 32128 13388 32180 13394
rect 32128 13330 32180 13336
rect 32232 13326 32260 14350
rect 32324 14006 32352 14350
rect 32312 14000 32364 14006
rect 32312 13942 32364 13948
rect 32324 13394 32352 13942
rect 32416 13938 32444 14894
rect 32496 14884 32548 14890
rect 32496 14826 32548 14832
rect 32508 14618 32536 14826
rect 32496 14612 32548 14618
rect 32496 14554 32548 14560
rect 32404 13932 32456 13938
rect 32404 13874 32456 13880
rect 32312 13388 32364 13394
rect 32312 13330 32364 13336
rect 32220 13320 32272 13326
rect 32220 13262 32272 13268
rect 32324 13274 32352 13330
rect 32324 13246 32536 13274
rect 32312 13184 32364 13190
rect 32312 13126 32364 13132
rect 31220 12406 31340 12434
rect 31404 12406 31524 12434
rect 30932 10668 30984 10674
rect 30932 10610 30984 10616
rect 30932 10532 30984 10538
rect 30932 10474 30984 10480
rect 30840 10464 30892 10470
rect 30944 10441 30972 10474
rect 30840 10406 30892 10412
rect 30930 10432 30986 10441
rect 30564 10134 30616 10140
rect 30668 10118 30788 10146
rect 30668 10062 30696 10118
rect 30852 10062 30880 10406
rect 30930 10367 30986 10376
rect 30656 10056 30708 10062
rect 30656 9998 30708 10004
rect 30840 10056 30892 10062
rect 30840 9998 30892 10004
rect 28908 8492 28960 8498
rect 28908 8434 28960 8440
rect 30472 8492 30524 8498
rect 30472 8434 30524 8440
rect 30668 8362 30696 9998
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 30760 8634 30788 8842
rect 30748 8628 30800 8634
rect 30748 8570 30800 8576
rect 30656 8356 30708 8362
rect 30656 8298 30708 8304
rect 30196 8288 30248 8294
rect 30196 8230 30248 8236
rect 30208 7818 30236 8230
rect 30668 7886 30696 8298
rect 30656 7880 30708 7886
rect 30656 7822 30708 7828
rect 30196 7812 30248 7818
rect 30196 7754 30248 7760
rect 29644 7744 29696 7750
rect 29644 7686 29696 7692
rect 29656 7410 29684 7686
rect 29644 7404 29696 7410
rect 29644 7346 29696 7352
rect 29828 7336 29880 7342
rect 29828 7278 29880 7284
rect 29644 7268 29696 7274
rect 29644 7210 29696 7216
rect 29460 4208 29512 4214
rect 29460 4150 29512 4156
rect 29472 3126 29500 4150
rect 29552 3528 29604 3534
rect 29552 3470 29604 3476
rect 29460 3120 29512 3126
rect 29460 3062 29512 3068
rect 29564 3058 29592 3470
rect 29552 3052 29604 3058
rect 29552 2994 29604 3000
rect 28724 1964 28776 1970
rect 28724 1906 28776 1912
rect 29656 800 29684 7210
rect 29840 7002 29868 7278
rect 29828 6996 29880 7002
rect 29828 6938 29880 6944
rect 30472 4616 30524 4622
rect 30472 4558 30524 4564
rect 30840 4616 30892 4622
rect 30840 4558 30892 4564
rect 30196 4140 30248 4146
rect 30196 4082 30248 4088
rect 29736 3936 29788 3942
rect 29736 3878 29788 3884
rect 29748 3058 29776 3878
rect 30208 3670 30236 4082
rect 30012 3664 30064 3670
rect 30012 3606 30064 3612
rect 30196 3664 30248 3670
rect 30196 3606 30248 3612
rect 29920 3392 29972 3398
rect 29920 3334 29972 3340
rect 29932 3126 29960 3334
rect 30024 3194 30052 3606
rect 30208 3534 30236 3606
rect 30196 3528 30248 3534
rect 30196 3470 30248 3476
rect 30288 3392 30340 3398
rect 30288 3334 30340 3340
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 29920 3120 29972 3126
rect 29920 3062 29972 3068
rect 29736 3052 29788 3058
rect 29736 2994 29788 3000
rect 30194 2952 30250 2961
rect 30194 2887 30250 2896
rect 30208 1442 30236 2887
rect 30300 2514 30328 3334
rect 30484 2582 30512 4558
rect 30852 3602 30880 4558
rect 31024 3936 31076 3942
rect 31024 3878 31076 3884
rect 31036 3602 31064 3878
rect 30840 3596 30892 3602
rect 30840 3538 30892 3544
rect 31024 3596 31076 3602
rect 31024 3538 31076 3544
rect 31220 2990 31248 12406
rect 31300 4140 31352 4146
rect 31404 4128 31432 12406
rect 31852 8424 31904 8430
rect 31852 8366 31904 8372
rect 31864 8090 31892 8366
rect 31852 8084 31904 8090
rect 31852 8026 31904 8032
rect 32324 6914 32352 13126
rect 32508 11694 32536 13246
rect 32496 11688 32548 11694
rect 32496 11630 32548 11636
rect 32600 9178 32628 18702
rect 32692 15858 32720 18822
rect 33520 17354 33548 22066
rect 33888 21554 33916 22374
rect 33968 22024 34020 22030
rect 33968 21966 34020 21972
rect 33876 21548 33928 21554
rect 33876 21490 33928 21496
rect 33980 21146 34008 21966
rect 33968 21140 34020 21146
rect 33968 21082 34020 21088
rect 33692 20936 33744 20942
rect 33692 20878 33744 20884
rect 33704 19854 33732 20878
rect 33968 20256 34020 20262
rect 33968 20198 34020 20204
rect 33980 19854 34008 20198
rect 33692 19848 33744 19854
rect 33692 19790 33744 19796
rect 33876 19848 33928 19854
rect 33876 19790 33928 19796
rect 33968 19848 34020 19854
rect 33968 19790 34020 19796
rect 33888 19718 33916 19790
rect 33876 19712 33928 19718
rect 33876 19654 33928 19660
rect 33520 17326 33824 17354
rect 33508 17196 33560 17202
rect 33508 17138 33560 17144
rect 33048 16992 33100 16998
rect 33048 16934 33100 16940
rect 33060 16658 33088 16934
rect 33520 16794 33548 17138
rect 33508 16788 33560 16794
rect 33508 16730 33560 16736
rect 33048 16652 33100 16658
rect 33048 16594 33100 16600
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 32692 15830 32812 15858
rect 32680 14272 32732 14278
rect 32680 14214 32732 14220
rect 32692 14006 32720 14214
rect 32680 14000 32732 14006
rect 32680 13942 32732 13948
rect 32784 13190 32812 15830
rect 32968 15638 32996 16526
rect 33060 16182 33088 16594
rect 33048 16176 33100 16182
rect 33048 16118 33100 16124
rect 32956 15632 33008 15638
rect 32956 15574 33008 15580
rect 33324 15496 33376 15502
rect 33324 15438 33376 15444
rect 33232 15020 33284 15026
rect 33232 14962 33284 14968
rect 33244 14346 33272 14962
rect 33336 14482 33364 15438
rect 33324 14476 33376 14482
rect 33324 14418 33376 14424
rect 33232 14340 33284 14346
rect 33232 14282 33284 14288
rect 33796 13938 33824 17326
rect 33888 15026 33916 19654
rect 33968 15496 34020 15502
rect 33968 15438 34020 15444
rect 33980 15162 34008 15438
rect 33968 15156 34020 15162
rect 33968 15098 34020 15104
rect 33876 15020 33928 15026
rect 33876 14962 33928 14968
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 32772 13184 32824 13190
rect 32772 13126 32824 13132
rect 32588 9172 32640 9178
rect 32588 9114 32640 9120
rect 32600 8498 32628 9114
rect 32588 8492 32640 8498
rect 32588 8434 32640 8440
rect 32324 6886 32444 6914
rect 31352 4100 31432 4128
rect 31300 4082 31352 4088
rect 31484 3936 31536 3942
rect 31484 3878 31536 3884
rect 32128 3936 32180 3942
rect 32128 3878 32180 3884
rect 31496 3126 31524 3878
rect 31576 3596 31628 3602
rect 31576 3538 31628 3544
rect 31484 3120 31536 3126
rect 31484 3062 31536 3068
rect 31208 2984 31260 2990
rect 31300 2984 31352 2990
rect 31208 2926 31260 2932
rect 31298 2952 31300 2961
rect 31352 2952 31354 2961
rect 31298 2887 31354 2896
rect 30472 2576 30524 2582
rect 30472 2518 30524 2524
rect 30288 2508 30340 2514
rect 30288 2450 30340 2456
rect 30932 2508 30984 2514
rect 30932 2450 30984 2456
rect 30208 1414 30328 1442
rect 30300 800 30328 1414
rect 30944 800 30972 2450
rect 31588 800 31616 3538
rect 32140 3058 32168 3878
rect 32416 3670 32444 6886
rect 33796 3738 33824 13874
rect 34072 6914 34100 28426
rect 34336 27600 34388 27606
rect 34336 27542 34388 27548
rect 34244 22636 34296 22642
rect 34244 22578 34296 22584
rect 34152 22500 34204 22506
rect 34152 22442 34204 22448
rect 34164 22234 34192 22442
rect 34152 22228 34204 22234
rect 34152 22170 34204 22176
rect 34164 22030 34192 22170
rect 34256 22166 34284 22578
rect 34244 22160 34296 22166
rect 34244 22102 34296 22108
rect 34152 22024 34204 22030
rect 34152 21966 34204 21972
rect 34244 20460 34296 20466
rect 34164 20420 34244 20448
rect 34164 12434 34192 20420
rect 34244 20402 34296 20408
rect 34164 12406 34284 12434
rect 33980 6886 34100 6914
rect 33784 3732 33836 3738
rect 33784 3674 33836 3680
rect 32404 3664 32456 3670
rect 32404 3606 32456 3612
rect 33980 3466 34008 6886
rect 33968 3460 34020 3466
rect 33968 3402 34020 3408
rect 34256 3194 34284 12406
rect 34244 3188 34296 3194
rect 34244 3130 34296 3136
rect 34348 3126 34376 27542
rect 34440 24750 34468 49302
rect 34612 48136 34664 48142
rect 34612 48078 34664 48084
rect 34624 47530 34652 48078
rect 34716 47598 34744 51326
rect 34794 51200 34850 51326
rect 35438 51200 35494 52000
rect 36082 51354 36138 52000
rect 36082 51326 36308 51354
rect 36082 51200 36138 51326
rect 34934 49532 35242 49552
rect 34934 49530 34940 49532
rect 34996 49530 35020 49532
rect 35076 49530 35100 49532
rect 35156 49530 35180 49532
rect 35236 49530 35242 49532
rect 34996 49478 34998 49530
rect 35178 49478 35180 49530
rect 34934 49476 34940 49478
rect 34996 49476 35020 49478
rect 35076 49476 35100 49478
rect 35156 49476 35180 49478
rect 35236 49476 35242 49478
rect 34934 49456 35242 49476
rect 34888 49224 34940 49230
rect 34888 49166 34940 49172
rect 36176 49224 36228 49230
rect 36176 49166 36228 49172
rect 34796 48816 34848 48822
rect 34796 48758 34848 48764
rect 34808 48346 34836 48758
rect 34900 48754 34928 49166
rect 34888 48748 34940 48754
rect 34888 48690 34940 48696
rect 34934 48444 35242 48464
rect 34934 48442 34940 48444
rect 34996 48442 35020 48444
rect 35076 48442 35100 48444
rect 35156 48442 35180 48444
rect 35236 48442 35242 48444
rect 34996 48390 34998 48442
rect 35178 48390 35180 48442
rect 34934 48388 34940 48390
rect 34996 48388 35020 48390
rect 35076 48388 35100 48390
rect 35156 48388 35180 48390
rect 35236 48388 35242 48390
rect 34934 48368 35242 48388
rect 34796 48340 34848 48346
rect 34796 48282 34848 48288
rect 36188 48210 36216 49166
rect 36280 48210 36308 51326
rect 36726 51200 36782 52000
rect 37370 51354 37426 52000
rect 38014 51354 38070 52000
rect 38658 51354 38714 52000
rect 37370 51326 37504 51354
rect 37370 51200 37426 51326
rect 36740 48822 36768 51200
rect 37004 49768 37056 49774
rect 37004 49710 37056 49716
rect 36728 48816 36780 48822
rect 36728 48758 36780 48764
rect 36636 48272 36688 48278
rect 36636 48214 36688 48220
rect 36176 48204 36228 48210
rect 36176 48146 36228 48152
rect 36268 48204 36320 48210
rect 36268 48146 36320 48152
rect 35900 48068 35952 48074
rect 35900 48010 35952 48016
rect 35912 47734 35940 48010
rect 35900 47728 35952 47734
rect 35900 47670 35952 47676
rect 35808 47660 35860 47666
rect 35808 47602 35860 47608
rect 34704 47592 34756 47598
rect 34704 47534 34756 47540
rect 34612 47524 34664 47530
rect 34612 47466 34664 47472
rect 34520 34536 34572 34542
rect 34520 34478 34572 34484
rect 34532 34202 34560 34478
rect 34520 34196 34572 34202
rect 34520 34138 34572 34144
rect 34520 29844 34572 29850
rect 34520 29786 34572 29792
rect 34532 29170 34560 29786
rect 34624 29730 34652 47466
rect 34934 47356 35242 47376
rect 34934 47354 34940 47356
rect 34996 47354 35020 47356
rect 35076 47354 35100 47356
rect 35156 47354 35180 47356
rect 35236 47354 35242 47356
rect 34996 47302 34998 47354
rect 35178 47302 35180 47354
rect 34934 47300 34940 47302
rect 34996 47300 35020 47302
rect 35076 47300 35100 47302
rect 35156 47300 35180 47302
rect 35236 47300 35242 47302
rect 34934 47280 35242 47300
rect 35820 47190 35848 47602
rect 35808 47184 35860 47190
rect 35808 47126 35860 47132
rect 34934 46268 35242 46288
rect 34934 46266 34940 46268
rect 34996 46266 35020 46268
rect 35076 46266 35100 46268
rect 35156 46266 35180 46268
rect 35236 46266 35242 46268
rect 34996 46214 34998 46266
rect 35178 46214 35180 46266
rect 34934 46212 34940 46214
rect 34996 46212 35020 46214
rect 35076 46212 35100 46214
rect 35156 46212 35180 46214
rect 35236 46212 35242 46214
rect 34934 46192 35242 46212
rect 34934 45180 35242 45200
rect 34934 45178 34940 45180
rect 34996 45178 35020 45180
rect 35076 45178 35100 45180
rect 35156 45178 35180 45180
rect 35236 45178 35242 45180
rect 34996 45126 34998 45178
rect 35178 45126 35180 45178
rect 34934 45124 34940 45126
rect 34996 45124 35020 45126
rect 35076 45124 35100 45126
rect 35156 45124 35180 45126
rect 35236 45124 35242 45126
rect 34934 45104 35242 45124
rect 36544 44328 36596 44334
rect 36544 44270 36596 44276
rect 34934 44092 35242 44112
rect 34934 44090 34940 44092
rect 34996 44090 35020 44092
rect 35076 44090 35100 44092
rect 35156 44090 35180 44092
rect 35236 44090 35242 44092
rect 34996 44038 34998 44090
rect 35178 44038 35180 44090
rect 34934 44036 34940 44038
rect 34996 44036 35020 44038
rect 35076 44036 35100 44038
rect 35156 44036 35180 44038
rect 35236 44036 35242 44038
rect 34934 44016 35242 44036
rect 34934 43004 35242 43024
rect 34934 43002 34940 43004
rect 34996 43002 35020 43004
rect 35076 43002 35100 43004
rect 35156 43002 35180 43004
rect 35236 43002 35242 43004
rect 34996 42950 34998 43002
rect 35178 42950 35180 43002
rect 34934 42948 34940 42950
rect 34996 42948 35020 42950
rect 35076 42948 35100 42950
rect 35156 42948 35180 42950
rect 35236 42948 35242 42950
rect 34934 42928 35242 42948
rect 34934 41916 35242 41936
rect 34934 41914 34940 41916
rect 34996 41914 35020 41916
rect 35076 41914 35100 41916
rect 35156 41914 35180 41916
rect 35236 41914 35242 41916
rect 34996 41862 34998 41914
rect 35178 41862 35180 41914
rect 34934 41860 34940 41862
rect 34996 41860 35020 41862
rect 35076 41860 35100 41862
rect 35156 41860 35180 41862
rect 35236 41860 35242 41862
rect 34934 41840 35242 41860
rect 34934 40828 35242 40848
rect 34934 40826 34940 40828
rect 34996 40826 35020 40828
rect 35076 40826 35100 40828
rect 35156 40826 35180 40828
rect 35236 40826 35242 40828
rect 34996 40774 34998 40826
rect 35178 40774 35180 40826
rect 34934 40772 34940 40774
rect 34996 40772 35020 40774
rect 35076 40772 35100 40774
rect 35156 40772 35180 40774
rect 35236 40772 35242 40774
rect 34934 40752 35242 40772
rect 34934 39740 35242 39760
rect 34934 39738 34940 39740
rect 34996 39738 35020 39740
rect 35076 39738 35100 39740
rect 35156 39738 35180 39740
rect 35236 39738 35242 39740
rect 34996 39686 34998 39738
rect 35178 39686 35180 39738
rect 34934 39684 34940 39686
rect 34996 39684 35020 39686
rect 35076 39684 35100 39686
rect 35156 39684 35180 39686
rect 35236 39684 35242 39686
rect 34934 39664 35242 39684
rect 34934 38652 35242 38672
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38576 35242 38596
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 35348 32836 35400 32842
rect 35348 32778 35400 32784
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 35360 32026 35388 32778
rect 35348 32020 35400 32026
rect 35348 31962 35400 31968
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 35440 30184 35492 30190
rect 35440 30126 35492 30132
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 34624 29702 34928 29730
rect 34612 29640 34664 29646
rect 34612 29582 34664 29588
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34624 28558 34652 29582
rect 34796 29504 34848 29510
rect 34796 29446 34848 29452
rect 34704 29096 34756 29102
rect 34704 29038 34756 29044
rect 34716 28762 34744 29038
rect 34704 28756 34756 28762
rect 34704 28698 34756 28704
rect 34612 28552 34664 28558
rect 34612 28494 34664 28500
rect 34624 27674 34652 28494
rect 34808 28150 34836 29446
rect 34900 29034 34928 29702
rect 34888 29028 34940 29034
rect 34888 28970 34940 28976
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 34796 28144 34848 28150
rect 34796 28086 34848 28092
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34612 27668 34664 27674
rect 34612 27610 34664 27616
rect 34704 27464 34756 27470
rect 34704 27406 34756 27412
rect 34716 27130 34744 27406
rect 34704 27124 34756 27130
rect 34704 27066 34756 27072
rect 34796 26988 34848 26994
rect 34796 26930 34848 26936
rect 34704 26920 34756 26926
rect 34704 26862 34756 26868
rect 34428 24744 34480 24750
rect 34428 24686 34480 24692
rect 34520 22432 34572 22438
rect 34520 22374 34572 22380
rect 34532 21962 34560 22374
rect 34612 22228 34664 22234
rect 34612 22170 34664 22176
rect 34520 21956 34572 21962
rect 34520 21898 34572 21904
rect 34428 20460 34480 20466
rect 34428 20402 34480 20408
rect 34440 19990 34468 20402
rect 34532 20398 34560 21898
rect 34624 20466 34652 22170
rect 34716 22094 34744 26862
rect 34808 26382 34836 26930
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34796 26376 34848 26382
rect 34796 26318 34848 26324
rect 35164 26240 35216 26246
rect 35164 26182 35216 26188
rect 35176 25906 35204 26182
rect 35164 25900 35216 25906
rect 35164 25842 35216 25848
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34796 25152 34848 25158
rect 34796 25094 34848 25100
rect 34808 24342 34836 25094
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34796 24336 34848 24342
rect 34796 24278 34848 24284
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 34716 22066 34836 22094
rect 34704 22024 34756 22030
rect 34704 21966 34756 21972
rect 34716 21622 34744 21966
rect 34704 21616 34756 21622
rect 34704 21558 34756 21564
rect 34716 20534 34744 21558
rect 34704 20528 34756 20534
rect 34704 20470 34756 20476
rect 34612 20460 34664 20466
rect 34612 20402 34664 20408
rect 34520 20392 34572 20398
rect 34520 20334 34572 20340
rect 34428 19984 34480 19990
rect 34428 19926 34480 19932
rect 34716 19922 34744 20470
rect 34704 19916 34756 19922
rect 34704 19858 34756 19864
rect 34808 4690 34836 22066
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 34796 4684 34848 4690
rect 34796 4626 34848 4632
rect 34520 4548 34572 4554
rect 34520 4490 34572 4496
rect 34336 3120 34388 3126
rect 34336 3062 34388 3068
rect 32128 3052 32180 3058
rect 32128 2994 32180 3000
rect 34532 2990 34560 4490
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33508 2984 33560 2990
rect 33508 2926 33560 2932
rect 34520 2984 34572 2990
rect 34520 2926 34572 2932
rect 32220 2916 32272 2922
rect 32220 2858 32272 2864
rect 32232 800 32260 2858
rect 33140 2576 33192 2582
rect 33140 2518 33192 2524
rect 32864 2440 32916 2446
rect 32864 2382 32916 2388
rect 32876 800 32904 2382
rect 33152 2038 33180 2518
rect 33140 2032 33192 2038
rect 33140 1974 33192 1980
rect 33520 800 33548 2926
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 35360 2582 35388 5578
rect 35452 4826 35480 30126
rect 35532 30116 35584 30122
rect 35532 30058 35584 30064
rect 35544 29714 35572 30058
rect 35532 29708 35584 29714
rect 35532 29650 35584 29656
rect 35716 29572 35768 29578
rect 35716 29514 35768 29520
rect 35728 29306 35756 29514
rect 35716 29300 35768 29306
rect 35716 29242 35768 29248
rect 36360 29096 36412 29102
rect 36360 29038 36412 29044
rect 35532 28552 35584 28558
rect 35532 28494 35584 28500
rect 35544 27946 35572 28494
rect 35716 28484 35768 28490
rect 35716 28426 35768 28432
rect 35728 28218 35756 28426
rect 35716 28212 35768 28218
rect 35716 28154 35768 28160
rect 35532 27940 35584 27946
rect 35532 27882 35584 27888
rect 35808 26988 35860 26994
rect 35808 26930 35860 26936
rect 35820 26246 35848 26930
rect 36268 26784 36320 26790
rect 36268 26726 36320 26732
rect 36280 26450 36308 26726
rect 36268 26444 36320 26450
rect 36268 26386 36320 26392
rect 35808 26240 35860 26246
rect 35808 26182 35860 26188
rect 35808 25832 35860 25838
rect 35808 25774 35860 25780
rect 35624 24608 35676 24614
rect 35624 24550 35676 24556
rect 35636 24342 35664 24550
rect 35624 24336 35676 24342
rect 35624 24278 35676 24284
rect 35440 4820 35492 4826
rect 35440 4762 35492 4768
rect 35820 3670 35848 25774
rect 36084 21888 36136 21894
rect 36084 21830 36136 21836
rect 36096 20942 36124 21830
rect 36084 20936 36136 20942
rect 36084 20878 36136 20884
rect 36372 5166 36400 29038
rect 36452 28008 36504 28014
rect 36452 27950 36504 27956
rect 36464 12442 36492 27950
rect 36556 24274 36584 44270
rect 36544 24268 36596 24274
rect 36544 24210 36596 24216
rect 36648 22234 36676 48214
rect 37016 32978 37044 49710
rect 37004 32972 37056 32978
rect 37004 32914 37056 32920
rect 37280 31816 37332 31822
rect 37280 31758 37332 31764
rect 37292 29170 37320 31758
rect 37476 29238 37504 51326
rect 38014 51326 38240 51354
rect 38014 51200 38070 51326
rect 38212 49230 38240 51326
rect 38658 51326 38884 51354
rect 38658 51200 38714 51326
rect 38200 49224 38252 49230
rect 38200 49166 38252 49172
rect 38016 49088 38068 49094
rect 38016 49030 38068 49036
rect 37464 29232 37516 29238
rect 37464 29174 37516 29180
rect 37280 29164 37332 29170
rect 37280 29106 37332 29112
rect 37188 28620 37240 28626
rect 37188 28562 37240 28568
rect 37096 27532 37148 27538
rect 37096 27474 37148 27480
rect 36636 22228 36688 22234
rect 36636 22170 36688 22176
rect 36544 21888 36596 21894
rect 36544 21830 36596 21836
rect 36556 21078 36584 21830
rect 36544 21072 36596 21078
rect 36544 21014 36596 21020
rect 36636 12776 36688 12782
rect 36636 12718 36688 12724
rect 36452 12436 36504 12442
rect 36452 12378 36504 12384
rect 36648 11762 36676 12718
rect 36636 11756 36688 11762
rect 36636 11698 36688 11704
rect 37108 6866 37136 27474
rect 37096 6860 37148 6866
rect 37096 6802 37148 6808
rect 37200 6730 37228 28562
rect 37292 28082 37320 29106
rect 37280 28076 37332 28082
rect 37280 28018 37332 28024
rect 37292 26994 37320 28018
rect 37372 27396 37424 27402
rect 37372 27338 37424 27344
rect 37384 27130 37412 27338
rect 37372 27124 37424 27130
rect 37372 27066 37424 27072
rect 37280 26988 37332 26994
rect 37280 26930 37332 26936
rect 38028 24818 38056 49030
rect 38856 31210 38884 51326
rect 39302 51200 39358 52000
rect 39946 51200 40002 52000
rect 40590 51354 40646 52000
rect 41234 51354 41290 52000
rect 41878 51354 41934 52000
rect 40590 51326 40816 51354
rect 40590 51200 40646 51326
rect 39316 46986 39344 51200
rect 39396 48680 39448 48686
rect 39960 48668 39988 51200
rect 40788 49162 40816 51326
rect 41234 51326 41368 51354
rect 41234 51200 41290 51326
rect 40776 49156 40828 49162
rect 40776 49098 40828 49104
rect 40868 49088 40920 49094
rect 40868 49030 40920 49036
rect 40040 48680 40092 48686
rect 39960 48640 40040 48668
rect 39396 48622 39448 48628
rect 40040 48622 40092 48628
rect 39408 48346 39436 48622
rect 39396 48340 39448 48346
rect 39396 48282 39448 48288
rect 39304 46980 39356 46986
rect 39304 46922 39356 46928
rect 40880 33590 40908 49030
rect 40868 33584 40920 33590
rect 40868 33526 40920 33532
rect 38844 31204 38896 31210
rect 38844 31146 38896 31152
rect 40132 30728 40184 30734
rect 40132 30670 40184 30676
rect 38476 25424 38528 25430
rect 38476 25366 38528 25372
rect 38106 24848 38162 24857
rect 38016 24812 38068 24818
rect 38106 24783 38162 24792
rect 38292 24812 38344 24818
rect 38016 24754 38068 24760
rect 38120 24750 38148 24783
rect 38292 24754 38344 24760
rect 38108 24744 38160 24750
rect 38108 24686 38160 24692
rect 38108 24608 38160 24614
rect 38108 24550 38160 24556
rect 37832 12708 37884 12714
rect 37832 12650 37884 12656
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 36360 5160 36412 5166
rect 36360 5102 36412 5108
rect 37372 4684 37424 4690
rect 37372 4626 37424 4632
rect 36268 3936 36320 3942
rect 36268 3878 36320 3884
rect 35808 3664 35860 3670
rect 35808 3606 35860 3612
rect 36280 3602 36308 3878
rect 36268 3596 36320 3602
rect 36268 3538 36320 3544
rect 36728 3596 36780 3602
rect 36728 3538 36780 3544
rect 36084 3528 36136 3534
rect 36084 3470 36136 3476
rect 36096 3058 36124 3470
rect 36084 3052 36136 3058
rect 36084 2994 36136 3000
rect 35072 2576 35124 2582
rect 35070 2544 35072 2553
rect 35348 2576 35400 2582
rect 35124 2544 35126 2553
rect 35348 2518 35400 2524
rect 35070 2479 35126 2488
rect 34796 2440 34848 2446
rect 34796 2382 34848 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 34152 2372 34204 2378
rect 34152 2314 34204 2320
rect 34164 800 34192 2314
rect 34808 800 34836 2382
rect 36096 800 36124 2382
rect 36740 800 36768 3538
rect 37384 800 37412 4626
rect 37844 4146 37872 12650
rect 37832 4140 37884 4146
rect 37832 4082 37884 4088
rect 38016 2984 38068 2990
rect 38016 2926 38068 2932
rect 38028 800 38056 2926
rect 38120 2378 38148 24550
rect 38304 8838 38332 24754
rect 38488 24614 38516 25366
rect 40144 25226 40172 30670
rect 40132 25220 40184 25226
rect 40132 25162 40184 25168
rect 40040 24744 40092 24750
rect 40040 24686 40092 24692
rect 38660 24676 38712 24682
rect 38660 24618 38712 24624
rect 38476 24608 38528 24614
rect 38476 24550 38528 24556
rect 38672 24410 38700 24618
rect 38660 24404 38712 24410
rect 38660 24346 38712 24352
rect 40052 24138 40080 24686
rect 40144 24206 40172 25162
rect 40224 24744 40276 24750
rect 40224 24686 40276 24692
rect 41236 24744 41288 24750
rect 41340 24732 41368 51326
rect 41708 51326 41934 51354
rect 41708 49162 41736 51326
rect 41878 51200 41934 51326
rect 42522 51200 42578 52000
rect 43166 51200 43222 52000
rect 43810 51354 43866 52000
rect 43810 51326 43944 51354
rect 43810 51200 43866 51326
rect 41696 49156 41748 49162
rect 41696 49098 41748 49104
rect 41788 49156 41840 49162
rect 41788 49098 41840 49104
rect 41604 49088 41656 49094
rect 41604 49030 41656 49036
rect 41420 48680 41472 48686
rect 41420 48622 41472 48628
rect 41432 47666 41460 48622
rect 41420 47660 41472 47666
rect 41420 47602 41472 47608
rect 41512 46980 41564 46986
rect 41512 46922 41564 46928
rect 41524 30938 41552 46922
rect 41512 30932 41564 30938
rect 41512 30874 41564 30880
rect 41288 24704 41368 24732
rect 41236 24686 41288 24692
rect 40236 24410 40264 24686
rect 40224 24404 40276 24410
rect 40224 24346 40276 24352
rect 40132 24200 40184 24206
rect 40132 24142 40184 24148
rect 40040 24132 40092 24138
rect 40040 24074 40092 24080
rect 41616 20330 41644 49030
rect 41800 48890 41828 49098
rect 41788 48884 41840 48890
rect 41788 48826 41840 48832
rect 41696 48748 41748 48754
rect 41696 48690 41748 48696
rect 41708 47802 41736 48690
rect 42536 48210 42564 51200
rect 43180 49298 43208 51200
rect 43168 49292 43220 49298
rect 43168 49234 43220 49240
rect 43076 48680 43128 48686
rect 43076 48622 43128 48628
rect 42524 48204 42576 48210
rect 42524 48146 42576 48152
rect 41788 48068 41840 48074
rect 41788 48010 41840 48016
rect 41696 47796 41748 47802
rect 41696 47738 41748 47744
rect 41800 46986 41828 48010
rect 43088 47802 43116 48622
rect 43916 48142 43944 51326
rect 44454 51200 44510 52000
rect 45098 51200 45154 52000
rect 45742 51200 45798 52000
rect 46386 51200 46442 52000
rect 46570 51776 46626 51785
rect 46570 51711 46626 51720
rect 43996 49224 44048 49230
rect 43996 49166 44048 49172
rect 43904 48136 43956 48142
rect 43904 48078 43956 48084
rect 43076 47796 43128 47802
rect 43076 47738 43128 47744
rect 42708 47660 42760 47666
rect 42708 47602 42760 47608
rect 42340 47252 42392 47258
rect 42340 47194 42392 47200
rect 42352 46986 42380 47194
rect 42720 47054 42748 47602
rect 42800 47592 42852 47598
rect 42800 47534 42852 47540
rect 42708 47048 42760 47054
rect 42708 46990 42760 46996
rect 41788 46980 41840 46986
rect 41788 46922 41840 46928
rect 42340 46980 42392 46986
rect 42340 46922 42392 46928
rect 41604 20324 41656 20330
rect 41604 20266 41656 20272
rect 38292 8832 38344 8838
rect 38292 8774 38344 8780
rect 38660 6452 38712 6458
rect 38660 6394 38712 6400
rect 38568 3528 38620 3534
rect 38568 3470 38620 3476
rect 38580 3058 38608 3470
rect 38568 3052 38620 3058
rect 38568 2994 38620 3000
rect 38672 2582 38700 6394
rect 42064 4548 42116 4554
rect 42064 4490 42116 4496
rect 42076 4282 42104 4490
rect 42064 4276 42116 4282
rect 42064 4218 42116 4224
rect 42352 4146 42380 46922
rect 42720 46578 42748 46990
rect 42708 46572 42760 46578
rect 42708 46514 42760 46520
rect 42720 46170 42748 46514
rect 42812 46510 42840 47534
rect 43628 47116 43680 47122
rect 43628 47058 43680 47064
rect 42800 46504 42852 46510
rect 42800 46446 42852 46452
rect 42708 46164 42760 46170
rect 42708 46106 42760 46112
rect 43444 44260 43496 44266
rect 43444 44202 43496 44208
rect 43456 34678 43484 44202
rect 43640 40050 43668 47058
rect 44008 46170 44036 49166
rect 44088 49156 44140 49162
rect 44088 49098 44140 49104
rect 44100 46714 44128 49098
rect 44468 48142 44496 51200
rect 45112 49314 45140 51200
rect 45558 51096 45614 51105
rect 45558 51031 45614 51040
rect 45572 49774 45600 51031
rect 45560 49768 45612 49774
rect 45560 49710 45612 49716
rect 45112 49298 45232 49314
rect 45112 49292 45244 49298
rect 45112 49286 45192 49292
rect 45192 49234 45244 49240
rect 45756 48686 45784 51200
rect 44824 48680 44876 48686
rect 44824 48622 44876 48628
rect 45376 48680 45428 48686
rect 45376 48622 45428 48628
rect 45744 48680 45796 48686
rect 45744 48622 45796 48628
rect 44456 48136 44508 48142
rect 44456 48078 44508 48084
rect 44364 48000 44416 48006
rect 44364 47942 44416 47948
rect 44088 46708 44140 46714
rect 44088 46650 44140 46656
rect 44180 46504 44232 46510
rect 44180 46446 44232 46452
rect 43996 46164 44048 46170
rect 43996 46106 44048 46112
rect 44192 45490 44220 46446
rect 44376 45966 44404 47942
rect 44732 47116 44784 47122
rect 44732 47058 44784 47064
rect 44364 45960 44416 45966
rect 44364 45902 44416 45908
rect 44744 45490 44772 47058
rect 44836 46170 44864 48622
rect 44916 48000 44968 48006
rect 44916 47942 44968 47948
rect 44824 46164 44876 46170
rect 44824 46106 44876 46112
rect 44180 45484 44232 45490
rect 44180 45426 44232 45432
rect 44732 45484 44784 45490
rect 44732 45426 44784 45432
rect 43628 40044 43680 40050
rect 43628 39986 43680 39992
rect 43444 34672 43496 34678
rect 43444 34614 43496 34620
rect 42800 30796 42852 30802
rect 42800 30738 42852 30744
rect 42812 29714 42840 30738
rect 42800 29708 42852 29714
rect 42800 29650 42852 29656
rect 44824 26308 44876 26314
rect 44824 26250 44876 26256
rect 44836 16833 44864 26250
rect 44928 24614 44956 47942
rect 45100 47592 45152 47598
rect 45100 47534 45152 47540
rect 45284 47592 45336 47598
rect 45284 47534 45336 47540
rect 45008 47048 45060 47054
rect 45008 46990 45060 46996
rect 45020 46646 45048 46990
rect 45008 46640 45060 46646
rect 45008 46582 45060 46588
rect 45112 44402 45140 47534
rect 45296 47258 45324 47534
rect 45284 47252 45336 47258
rect 45284 47194 45336 47200
rect 45388 46170 45416 48622
rect 46480 48068 46532 48074
rect 46480 48010 46532 48016
rect 45560 47728 45612 47734
rect 45560 47670 45612 47676
rect 45376 46164 45428 46170
rect 45376 46106 45428 46112
rect 45192 45416 45244 45422
rect 45192 45358 45244 45364
rect 45204 45082 45232 45358
rect 45572 45082 45600 47670
rect 45652 47048 45704 47054
rect 45652 46990 45704 46996
rect 45192 45076 45244 45082
rect 45192 45018 45244 45024
rect 45560 45076 45612 45082
rect 45560 45018 45612 45024
rect 45558 44976 45614 44985
rect 45558 44911 45614 44920
rect 45100 44396 45152 44402
rect 45100 44338 45152 44344
rect 45572 44334 45600 44911
rect 45560 44328 45612 44334
rect 45560 44270 45612 44276
rect 45664 44282 45692 46990
rect 45836 46980 45888 46986
rect 45836 46922 45888 46928
rect 45744 46912 45796 46918
rect 45744 46854 45796 46860
rect 45756 46646 45784 46854
rect 45744 46640 45796 46646
rect 45744 46582 45796 46588
rect 45848 45082 45876 46922
rect 46492 46170 46520 48010
rect 46584 47598 46612 51711
rect 47030 51200 47086 52000
rect 47674 51354 47730 52000
rect 47674 51326 47808 51354
rect 47674 51200 47730 51326
rect 46846 50416 46902 50425
rect 46846 50351 46902 50360
rect 46754 49736 46810 49745
rect 46754 49671 46810 49680
rect 46664 48204 46716 48210
rect 46664 48146 46716 48152
rect 46572 47592 46624 47598
rect 46572 47534 46624 47540
rect 46572 47456 46624 47462
rect 46572 47398 46624 47404
rect 46480 46164 46532 46170
rect 46480 46106 46532 46112
rect 46296 45960 46348 45966
rect 46296 45902 46348 45908
rect 45836 45076 45888 45082
rect 45836 45018 45888 45024
rect 45928 44872 45980 44878
rect 45928 44814 45980 44820
rect 45664 44254 45876 44282
rect 45652 44192 45704 44198
rect 45652 44134 45704 44140
rect 45558 26616 45614 26625
rect 45558 26551 45614 26560
rect 45572 25974 45600 26551
rect 45560 25968 45612 25974
rect 45560 25910 45612 25916
rect 45664 24818 45692 44134
rect 45744 42288 45796 42294
rect 45744 42230 45796 42236
rect 45756 26518 45784 42230
rect 45848 29170 45876 44254
rect 45940 44198 45968 44814
rect 46308 44402 46336 45902
rect 46584 44402 46612 47398
rect 46296 44396 46348 44402
rect 46296 44338 46348 44344
rect 46572 44396 46624 44402
rect 46572 44338 46624 44344
rect 46018 44296 46074 44305
rect 46584 44282 46612 44338
rect 46018 44231 46020 44240
rect 46072 44231 46074 44240
rect 46400 44254 46612 44282
rect 46020 44202 46072 44208
rect 45928 44192 45980 44198
rect 45928 44134 45980 44140
rect 46296 39840 46348 39846
rect 46296 39782 46348 39788
rect 46308 39506 46336 39782
rect 46296 39500 46348 39506
rect 46296 39442 46348 39448
rect 46296 37256 46348 37262
rect 46296 37198 46348 37204
rect 46308 36786 46336 37198
rect 46400 36854 46428 44254
rect 46676 43926 46704 48146
rect 46768 47122 46796 49671
rect 46860 48210 46888 50351
rect 47780 49230 47808 51326
rect 48318 51200 48374 52000
rect 48962 51200 49018 52000
rect 49606 51200 49662 52000
rect 47768 49224 47820 49230
rect 47768 49166 47820 49172
rect 47308 49088 47360 49094
rect 47308 49030 47360 49036
rect 47766 49056 47822 49065
rect 47124 48544 47176 48550
rect 47124 48486 47176 48492
rect 47032 48272 47084 48278
rect 47032 48214 47084 48220
rect 46848 48204 46900 48210
rect 46848 48146 46900 48152
rect 46756 47116 46808 47122
rect 46756 47058 46808 47064
rect 46846 47016 46902 47025
rect 46846 46951 46902 46960
rect 46756 46028 46808 46034
rect 46756 45970 46808 45976
rect 46768 45234 46796 45970
rect 46860 45422 46888 46951
rect 47044 46646 47072 48214
rect 47032 46640 47084 46646
rect 47032 46582 47084 46588
rect 46848 45416 46900 45422
rect 46848 45358 46900 45364
rect 46768 45206 46888 45234
rect 46756 44940 46808 44946
rect 46756 44882 46808 44888
rect 46768 43994 46796 44882
rect 46756 43988 46808 43994
rect 46756 43930 46808 43936
rect 46664 43920 46716 43926
rect 46664 43862 46716 43868
rect 46480 42628 46532 42634
rect 46480 42570 46532 42576
rect 46492 42294 46520 42570
rect 46480 42288 46532 42294
rect 46480 42230 46532 42236
rect 46480 41540 46532 41546
rect 46480 41482 46532 41488
rect 46492 41274 46520 41482
rect 46860 41414 46888 45206
rect 46940 44804 46992 44810
rect 46940 44746 46992 44752
rect 46952 44538 46980 44746
rect 46940 44532 46992 44538
rect 46940 44474 46992 44480
rect 46940 43648 46992 43654
rect 46940 43590 46992 43596
rect 46676 41386 46888 41414
rect 46676 41290 46704 41386
rect 46480 41268 46532 41274
rect 46480 41210 46532 41216
rect 46584 41262 46704 41290
rect 46388 36848 46440 36854
rect 46388 36790 46440 36796
rect 46296 36780 46348 36786
rect 46296 36722 46348 36728
rect 46480 35012 46532 35018
rect 46480 34954 46532 34960
rect 46296 34400 46348 34406
rect 46296 34342 46348 34348
rect 45928 33516 45980 33522
rect 45928 33458 45980 33464
rect 45836 29164 45888 29170
rect 45836 29106 45888 29112
rect 45744 26512 45796 26518
rect 45744 26454 45796 26460
rect 45940 26450 45968 33458
rect 46308 32978 46336 34342
rect 46492 33658 46520 34954
rect 46480 33652 46532 33658
rect 46480 33594 46532 33600
rect 46584 33522 46612 41262
rect 46664 41132 46716 41138
rect 46664 41074 46716 41080
rect 46572 33516 46624 33522
rect 46572 33458 46624 33464
rect 46480 33312 46532 33318
rect 46480 33254 46532 33260
rect 46492 32978 46520 33254
rect 46296 32972 46348 32978
rect 46296 32914 46348 32920
rect 46480 32972 46532 32978
rect 46480 32914 46532 32920
rect 46584 26586 46612 33458
rect 46572 26580 46624 26586
rect 46572 26522 46624 26528
rect 45928 26444 45980 26450
rect 45928 26386 45980 26392
rect 46676 25838 46704 41074
rect 46952 38434 46980 43590
rect 47032 43104 47084 43110
rect 47032 43046 47084 43052
rect 47044 42770 47072 43046
rect 47032 42764 47084 42770
rect 47032 42706 47084 42712
rect 47032 38752 47084 38758
rect 47032 38694 47084 38700
rect 46860 38406 46980 38434
rect 47044 38418 47072 38694
rect 47032 38412 47084 38418
rect 46860 37890 46888 38406
rect 47032 38354 47084 38360
rect 46940 38276 46992 38282
rect 46940 38218 46992 38224
rect 46952 38010 46980 38218
rect 46940 38004 46992 38010
rect 46940 37946 46992 37952
rect 46860 37862 46980 37890
rect 46846 37496 46902 37505
rect 46846 37431 46902 37440
rect 46860 37330 46888 37431
rect 46848 37324 46900 37330
rect 46848 37266 46900 37272
rect 46848 29572 46900 29578
rect 46848 29514 46900 29520
rect 46860 29345 46888 29514
rect 46846 29336 46902 29345
rect 46846 29271 46902 29280
rect 46664 25832 46716 25838
rect 46664 25774 46716 25780
rect 45652 24812 45704 24818
rect 45652 24754 45704 24760
rect 44916 24608 44968 24614
rect 44916 24550 44968 24556
rect 46296 24608 46348 24614
rect 46296 24550 46348 24556
rect 46308 24274 46336 24550
rect 46296 24268 46348 24274
rect 46296 24210 46348 24216
rect 46952 22710 46980 37862
rect 47032 35148 47084 35154
rect 47032 35090 47084 35096
rect 47044 34474 47072 35090
rect 47032 34468 47084 34474
rect 47032 34410 47084 34416
rect 47032 28960 47084 28966
rect 47032 28902 47084 28908
rect 47044 28626 47072 28902
rect 47032 28620 47084 28626
rect 47032 28562 47084 28568
rect 47136 28506 47164 48486
rect 47216 45824 47268 45830
rect 47216 45766 47268 45772
rect 47228 42226 47256 45766
rect 47320 43450 47348 49030
rect 47766 48991 47822 49000
rect 47780 48822 47808 48991
rect 48332 48890 48360 51200
rect 48320 48884 48372 48890
rect 48320 48826 48372 48832
rect 47768 48816 47820 48822
rect 47768 48758 47820 48764
rect 47766 48376 47822 48385
rect 47766 48311 47822 48320
rect 47780 47734 47808 48311
rect 47768 47728 47820 47734
rect 47768 47670 47820 47676
rect 47584 47456 47636 47462
rect 47584 47398 47636 47404
rect 47492 44396 47544 44402
rect 47492 44338 47544 44344
rect 47504 43722 47532 44338
rect 47492 43716 47544 43722
rect 47492 43658 47544 43664
rect 47308 43444 47360 43450
rect 47308 43386 47360 43392
rect 47216 42220 47268 42226
rect 47216 42162 47268 42168
rect 47306 40896 47362 40905
rect 47306 40831 47362 40840
rect 47320 40594 47348 40831
rect 47308 40588 47360 40594
rect 47308 40530 47360 40536
rect 47400 40520 47452 40526
rect 47400 40462 47452 40468
rect 47308 37868 47360 37874
rect 47308 37810 47360 37816
rect 47216 35488 47268 35494
rect 47216 35430 47268 35436
rect 47228 34134 47256 35430
rect 47320 34610 47348 37810
rect 47308 34604 47360 34610
rect 47308 34546 47360 34552
rect 47216 34128 47268 34134
rect 47216 34070 47268 34076
rect 47320 33946 47348 34546
rect 47228 33918 47348 33946
rect 47228 29458 47256 33918
rect 47306 30016 47362 30025
rect 47306 29951 47362 29960
rect 47320 29646 47348 29951
rect 47308 29640 47360 29646
rect 47308 29582 47360 29588
rect 47228 29430 47348 29458
rect 47216 29164 47268 29170
rect 47216 29106 47268 29112
rect 47044 28478 47164 28506
rect 46940 22704 46992 22710
rect 46940 22646 46992 22652
rect 47044 20058 47072 28478
rect 47228 26234 47256 29106
rect 47320 27606 47348 29430
rect 47308 27600 47360 27606
rect 47308 27542 47360 27548
rect 47308 27464 47360 27470
rect 47308 27406 47360 27412
rect 47136 26206 47256 26234
rect 47136 25498 47164 26206
rect 47124 25492 47176 25498
rect 47124 25434 47176 25440
rect 47216 24812 47268 24818
rect 47216 24754 47268 24760
rect 47032 20052 47084 20058
rect 47032 19994 47084 20000
rect 46756 19780 46808 19786
rect 46756 19722 46808 19728
rect 46768 19514 46796 19722
rect 46756 19508 46808 19514
rect 46756 19450 46808 19456
rect 46204 18760 46256 18766
rect 46204 18702 46256 18708
rect 45650 17776 45706 17785
rect 45650 17711 45706 17720
rect 45664 16833 45692 17711
rect 44822 16824 44878 16833
rect 44822 16759 44878 16768
rect 45650 16824 45706 16833
rect 45650 16759 45706 16768
rect 45560 12436 45612 12442
rect 45560 12378 45612 12384
rect 45572 12345 45600 12378
rect 45558 12336 45614 12345
rect 45558 12271 45614 12280
rect 42432 9988 42484 9994
rect 42432 9930 42484 9936
rect 42444 4146 42472 9930
rect 45744 7404 45796 7410
rect 45744 7346 45796 7352
rect 45558 6896 45614 6905
rect 45558 6831 45614 6840
rect 45652 6860 45704 6866
rect 45572 6730 45600 6831
rect 45652 6802 45704 6808
rect 45560 6724 45612 6730
rect 45560 6666 45612 6672
rect 45664 6225 45692 6802
rect 45650 6216 45706 6225
rect 45650 6151 45706 6160
rect 45560 4820 45612 4826
rect 45560 4762 45612 4768
rect 43076 4684 43128 4690
rect 43076 4626 43128 4632
rect 43260 4684 43312 4690
rect 43260 4626 43312 4632
rect 42340 4140 42392 4146
rect 42340 4082 42392 4088
rect 42432 4140 42484 4146
rect 42432 4082 42484 4088
rect 38752 3936 38804 3942
rect 38752 3878 38804 3884
rect 40776 3936 40828 3942
rect 40776 3878 40828 3884
rect 42432 3936 42484 3942
rect 42432 3878 42484 3884
rect 38764 2990 38792 3878
rect 40788 3602 40816 3878
rect 40776 3596 40828 3602
rect 40776 3538 40828 3544
rect 41236 3596 41288 3602
rect 41236 3538 41288 3544
rect 38752 2984 38804 2990
rect 38752 2926 38804 2932
rect 39948 2984 40000 2990
rect 39948 2926 40000 2932
rect 38660 2576 38712 2582
rect 38660 2518 38712 2524
rect 38660 2440 38712 2446
rect 38660 2382 38712 2388
rect 38108 2372 38160 2378
rect 38108 2314 38160 2320
rect 38672 800 38700 2382
rect 39960 800 39988 2926
rect 41248 800 41276 3538
rect 42444 3058 42472 3878
rect 43088 3738 43116 4626
rect 43076 3732 43128 3738
rect 43076 3674 43128 3680
rect 43272 3398 43300 4626
rect 44732 4616 44784 4622
rect 44732 4558 44784 4564
rect 43996 4140 44048 4146
rect 43996 4082 44048 4088
rect 43812 4072 43864 4078
rect 43812 4014 43864 4020
rect 43824 3738 43852 4014
rect 44008 3738 44036 4082
rect 44456 4072 44508 4078
rect 44456 4014 44508 4020
rect 43812 3732 43864 3738
rect 43812 3674 43864 3680
rect 43996 3732 44048 3738
rect 43996 3674 44048 3680
rect 42524 3392 42576 3398
rect 42524 3334 42576 3340
rect 43260 3392 43312 3398
rect 43260 3334 43312 3340
rect 42432 3052 42484 3058
rect 42432 2994 42484 3000
rect 41880 2848 41932 2854
rect 41880 2790 41932 2796
rect 41892 800 41920 2790
rect 42536 800 42564 3334
rect 42708 2984 42760 2990
rect 42708 2926 42760 2932
rect 42720 2854 42748 2926
rect 42708 2848 42760 2854
rect 42708 2790 42760 2796
rect 43168 2372 43220 2378
rect 43168 2314 43220 2320
rect 43180 800 43208 2314
rect 44468 800 44496 4014
rect 44744 3058 44772 4558
rect 45468 4140 45520 4146
rect 45468 4082 45520 4088
rect 44824 4004 44876 4010
rect 44824 3946 44876 3952
rect 44836 3466 44864 3946
rect 45480 3670 45508 4082
rect 45468 3664 45520 3670
rect 45468 3606 45520 3612
rect 45572 3505 45600 4762
rect 45756 3942 45784 7346
rect 45836 4616 45888 4622
rect 45836 4558 45888 4564
rect 45744 3936 45796 3942
rect 45744 3878 45796 3884
rect 45558 3496 45614 3505
rect 44824 3460 44876 3466
rect 45558 3431 45614 3440
rect 44824 3402 44876 3408
rect 44916 3392 44968 3398
rect 44916 3334 44968 3340
rect 44928 3126 44956 3334
rect 44916 3120 44968 3126
rect 44916 3062 44968 3068
rect 44732 3052 44784 3058
rect 44732 2994 44784 3000
rect 45100 2984 45152 2990
rect 45100 2926 45152 2932
rect 45112 800 45140 2926
rect 45848 2514 45876 4558
rect 46216 4185 46244 18702
rect 46296 17672 46348 17678
rect 46296 17614 46348 17620
rect 46308 16658 46336 17614
rect 46388 17264 46440 17270
rect 46388 17206 46440 17212
rect 46296 16652 46348 16658
rect 46296 16594 46348 16600
rect 46296 11552 46348 11558
rect 46296 11494 46348 11500
rect 46308 11218 46336 11494
rect 46296 11212 46348 11218
rect 46296 11154 46348 11160
rect 46400 9625 46428 17206
rect 47228 17202 47256 24754
rect 47320 23798 47348 27406
rect 47308 23792 47360 23798
rect 47308 23734 47360 23740
rect 47412 22098 47440 40462
rect 47492 40044 47544 40050
rect 47492 39986 47544 39992
rect 47504 32178 47532 39986
rect 47596 32314 47624 47398
rect 48976 47054 49004 51200
rect 49620 48278 49648 51200
rect 49608 48272 49660 48278
rect 49608 48214 49660 48220
rect 47952 47048 48004 47054
rect 47952 46990 48004 46996
rect 48964 47048 49016 47054
rect 48964 46990 49016 46996
rect 47964 46646 47992 46990
rect 47952 46640 48004 46646
rect 47952 46582 48004 46588
rect 47768 46368 47820 46374
rect 47768 46310 47820 46316
rect 48134 46336 48190 46345
rect 47676 45892 47728 45898
rect 47676 45834 47728 45840
rect 47688 45558 47716 45834
rect 47676 45552 47728 45558
rect 47676 45494 47728 45500
rect 47676 45348 47728 45354
rect 47676 45290 47728 45296
rect 47688 44538 47716 45290
rect 47676 44532 47728 44538
rect 47676 44474 47728 44480
rect 47676 41676 47728 41682
rect 47676 41618 47728 41624
rect 47688 41138 47716 41618
rect 47676 41132 47728 41138
rect 47676 41074 47728 41080
rect 47676 39840 47728 39846
rect 47676 39782 47728 39788
rect 47688 39506 47716 39782
rect 47676 39500 47728 39506
rect 47676 39442 47728 39448
rect 47676 37188 47728 37194
rect 47676 37130 47728 37136
rect 47688 36922 47716 37130
rect 47676 36916 47728 36922
rect 47676 36858 47728 36864
rect 47676 34400 47728 34406
rect 47676 34342 47728 34348
rect 47688 34066 47716 34342
rect 47676 34060 47728 34066
rect 47676 34002 47728 34008
rect 47596 32286 47716 32314
rect 47504 32150 47624 32178
rect 47490 32056 47546 32065
rect 47490 31991 47546 32000
rect 47504 31822 47532 31991
rect 47492 31816 47544 31822
rect 47492 31758 47544 31764
rect 47596 31090 47624 32150
rect 47504 31062 47624 31090
rect 47400 22092 47452 22098
rect 47400 22034 47452 22040
rect 47306 19136 47362 19145
rect 47306 19071 47362 19080
rect 47320 18834 47348 19071
rect 47308 18828 47360 18834
rect 47308 18770 47360 18776
rect 47216 17196 47268 17202
rect 47216 17138 47268 17144
rect 47032 16992 47084 16998
rect 47032 16934 47084 16940
rect 46480 15904 46532 15910
rect 46480 15846 46532 15852
rect 46492 15570 46520 15846
rect 47044 15638 47072 16934
rect 47228 16114 47256 17138
rect 47216 16108 47268 16114
rect 47216 16050 47268 16056
rect 47032 15632 47084 15638
rect 47032 15574 47084 15580
rect 46480 15564 46532 15570
rect 46480 15506 46532 15512
rect 46846 15056 46902 15065
rect 46846 14991 46848 15000
rect 46900 14991 46902 15000
rect 46848 14962 46900 14968
rect 46848 14340 46900 14346
rect 46848 14282 46900 14288
rect 46860 14074 46888 14282
rect 46848 14068 46900 14074
rect 46848 14010 46900 14016
rect 46846 13016 46902 13025
rect 46846 12951 46902 12960
rect 46860 12782 46888 12951
rect 46848 12776 46900 12782
rect 46848 12718 46900 12724
rect 46940 11076 46992 11082
rect 46940 11018 46992 11024
rect 46952 10810 46980 11018
rect 46940 10804 46992 10810
rect 46940 10746 46992 10752
rect 46848 10668 46900 10674
rect 46848 10610 46900 10616
rect 46860 9994 46888 10610
rect 46848 9988 46900 9994
rect 46848 9930 46900 9936
rect 46386 9616 46442 9625
rect 46386 9551 46442 9560
rect 46480 7200 46532 7206
rect 46480 7142 46532 7148
rect 46492 6866 46520 7142
rect 46480 6860 46532 6866
rect 46480 6802 46532 6808
rect 46848 5228 46900 5234
rect 46848 5170 46900 5176
rect 46756 4208 46808 4214
rect 46202 4176 46258 4185
rect 46756 4150 46808 4156
rect 46202 4111 46258 4120
rect 46204 3936 46256 3942
rect 46204 3878 46256 3884
rect 46216 3602 46244 3878
rect 46204 3596 46256 3602
rect 46204 3538 46256 3544
rect 46388 3596 46440 3602
rect 46388 3538 46440 3544
rect 45836 2508 45888 2514
rect 45836 2450 45888 2456
rect 45744 2304 45796 2310
rect 45744 2246 45796 2252
rect 45756 800 45784 2246
rect 46400 800 46428 3538
rect 11256 734 11560 762
rect 11610 0 11666 800
rect 12254 0 12310 800
rect 12898 0 12954 800
rect 13542 0 13598 800
rect 14186 0 14242 800
rect 14830 0 14886 800
rect 15474 0 15530 800
rect 16118 0 16174 800
rect 16762 0 16818 800
rect 17406 0 17462 800
rect 18050 0 18106 800
rect 18694 0 18750 800
rect 19338 0 19394 800
rect 19982 0 20038 800
rect 20626 0 20682 800
rect 21270 0 21326 800
rect 21914 0 21970 800
rect 22558 0 22614 800
rect 23202 0 23258 800
rect 23846 0 23902 800
rect 24490 0 24546 800
rect 25134 0 25190 800
rect 25778 0 25834 800
rect 26422 0 26478 800
rect 27066 0 27122 800
rect 27710 0 27766 800
rect 28354 0 28410 800
rect 28998 0 29054 800
rect 29642 0 29698 800
rect 30286 0 30342 800
rect 30930 0 30986 800
rect 31574 0 31630 800
rect 32218 0 32274 800
rect 32862 0 32918 800
rect 33506 0 33562 800
rect 34150 0 34206 800
rect 34794 0 34850 800
rect 35438 0 35494 800
rect 36082 0 36138 800
rect 36726 0 36782 800
rect 37370 0 37426 800
rect 38014 0 38070 800
rect 38658 0 38714 800
rect 39946 0 40002 800
rect 40590 0 40646 800
rect 41234 0 41290 800
rect 41878 0 41934 800
rect 42522 0 42578 800
rect 43166 0 43222 800
rect 43810 0 43866 800
rect 44454 0 44510 800
rect 45098 0 45154 800
rect 45742 0 45798 800
rect 46386 0 46442 800
rect 46768 105 46796 4150
rect 46860 4010 46888 5170
rect 47032 5160 47084 5166
rect 47032 5102 47084 5108
rect 46940 5024 46992 5030
rect 46940 4966 46992 4972
rect 46848 4004 46900 4010
rect 46848 3946 46900 3952
rect 46848 2644 46900 2650
rect 46848 2586 46900 2592
rect 46860 1465 46888 2586
rect 46952 2378 46980 4966
rect 46940 2372 46992 2378
rect 46940 2314 46992 2320
rect 46846 1456 46902 1465
rect 46846 1391 46902 1400
rect 47044 800 47072 5102
rect 47228 3466 47256 16050
rect 47400 5704 47452 5710
rect 47400 5646 47452 5652
rect 47412 4758 47440 5646
rect 47504 5234 47532 31062
rect 47688 30954 47716 32286
rect 47596 30926 47716 30954
rect 47596 23769 47624 30926
rect 47676 28960 47728 28966
rect 47676 28902 47728 28908
rect 47688 28490 47716 28902
rect 47676 28484 47728 28490
rect 47676 28426 47728 28432
rect 47676 28212 47728 28218
rect 47676 28154 47728 28160
rect 47688 27470 47716 28154
rect 47676 27464 47728 27470
rect 47676 27406 47728 27412
rect 47676 24608 47728 24614
rect 47676 24550 47728 24556
rect 47688 24274 47716 24550
rect 47676 24268 47728 24274
rect 47676 24210 47728 24216
rect 47582 23760 47638 23769
rect 47582 23695 47638 23704
rect 47584 22432 47636 22438
rect 47584 22374 47636 22380
rect 47596 22030 47624 22374
rect 47780 22234 47808 46310
rect 48134 46271 48190 46280
rect 48148 46034 48176 46271
rect 48136 46028 48188 46034
rect 48136 45970 48188 45976
rect 48134 45656 48190 45665
rect 48134 45591 48190 45600
rect 48148 44946 48176 45591
rect 48136 44940 48188 44946
rect 48136 44882 48188 44888
rect 47860 43784 47912 43790
rect 47860 43726 47912 43732
rect 47872 42945 47900 43726
rect 48228 43716 48280 43722
rect 48228 43658 48280 43664
rect 48134 43616 48190 43625
rect 48134 43551 48190 43560
rect 47952 43308 48004 43314
rect 47952 43250 48004 43256
rect 47858 42936 47914 42945
rect 47858 42871 47914 42880
rect 47964 42265 47992 43250
rect 48044 43104 48096 43110
rect 48044 43046 48096 43052
rect 47950 42256 48006 42265
rect 47860 42220 47912 42226
rect 47950 42191 48006 42200
rect 47860 42162 47912 42168
rect 47872 38706 47900 42162
rect 48056 41750 48084 43046
rect 48148 42770 48176 43551
rect 48136 42764 48188 42770
rect 48136 42706 48188 42712
rect 48044 41744 48096 41750
rect 48044 41686 48096 41692
rect 48134 41576 48190 41585
rect 48134 41511 48136 41520
rect 48188 41511 48190 41520
rect 48136 41482 48188 41488
rect 48134 40216 48190 40225
rect 48134 40151 48190 40160
rect 48044 39636 48096 39642
rect 48044 39578 48096 39584
rect 48056 39098 48084 39578
rect 48148 39506 48176 40151
rect 48240 39658 48268 43658
rect 48240 39630 48360 39658
rect 48226 39536 48282 39545
rect 48136 39500 48188 39506
rect 48226 39471 48282 39480
rect 48136 39442 48188 39448
rect 48044 39092 48096 39098
rect 48044 39034 48096 39040
rect 47952 38956 48004 38962
rect 47952 38898 48004 38904
rect 47964 38865 47992 38898
rect 47950 38856 48006 38865
rect 47950 38791 48006 38800
rect 47872 38678 47992 38706
rect 47858 38176 47914 38185
rect 47858 38111 47914 38120
rect 47872 37874 47900 38111
rect 47860 37868 47912 37874
rect 47860 37810 47912 37816
rect 47860 36168 47912 36174
rect 47858 36136 47860 36145
rect 47912 36136 47914 36145
rect 47858 36071 47914 36080
rect 47964 35894 47992 38678
rect 48240 38418 48268 39471
rect 48228 38412 48280 38418
rect 48228 38354 48280 38360
rect 48332 38298 48360 39630
rect 48240 38270 48360 38298
rect 48044 37664 48096 37670
rect 48044 37606 48096 37612
rect 47872 35866 47992 35894
rect 47872 31890 47900 35866
rect 48056 34218 48084 37606
rect 48136 37188 48188 37194
rect 48136 37130 48188 37136
rect 48148 36825 48176 37130
rect 48134 36816 48190 36825
rect 48134 36751 48190 36760
rect 48136 36032 48188 36038
rect 48136 35974 48188 35980
rect 48148 35578 48176 35974
rect 48240 35698 48268 38270
rect 48228 35692 48280 35698
rect 48228 35634 48280 35640
rect 48148 35550 48360 35578
rect 48228 35488 48280 35494
rect 48134 35456 48190 35465
rect 48228 35430 48280 35436
rect 48134 35391 48190 35400
rect 48148 35154 48176 35391
rect 48136 35148 48188 35154
rect 48136 35090 48188 35096
rect 48134 34776 48190 34785
rect 48134 34711 48190 34720
rect 47964 34190 48084 34218
rect 47964 33862 47992 34190
rect 48042 34096 48098 34105
rect 48148 34066 48176 34711
rect 48042 34031 48098 34040
rect 48136 34060 48188 34066
rect 47952 33856 48004 33862
rect 47952 33798 48004 33804
rect 47952 33516 48004 33522
rect 47952 33458 48004 33464
rect 47964 33425 47992 33458
rect 47950 33416 48006 33425
rect 47950 33351 48006 33360
rect 47952 33312 48004 33318
rect 47952 33254 48004 33260
rect 47860 31884 47912 31890
rect 47860 31826 47912 31832
rect 47964 31498 47992 33254
rect 48056 32978 48084 34031
rect 48136 34002 48188 34008
rect 48136 33856 48188 33862
rect 48136 33798 48188 33804
rect 48044 32972 48096 32978
rect 48044 32914 48096 32920
rect 47872 31470 47992 31498
rect 47872 28218 47900 31470
rect 47950 31376 48006 31385
rect 47950 31311 47952 31320
rect 48004 31311 48006 31320
rect 47952 31282 48004 31288
rect 48148 28778 48176 33798
rect 47964 28750 48176 28778
rect 47860 28212 47912 28218
rect 47860 28154 47912 28160
rect 47860 28076 47912 28082
rect 47860 28018 47912 28024
rect 47872 27985 47900 28018
rect 47858 27976 47914 27985
rect 47858 27911 47914 27920
rect 47964 27826 47992 28750
rect 48134 28656 48190 28665
rect 48134 28591 48136 28600
rect 48188 28591 48190 28600
rect 48136 28562 48188 28568
rect 47872 27798 47992 27826
rect 48044 27872 48096 27878
rect 48044 27814 48096 27820
rect 47872 25378 47900 27798
rect 47952 26308 48004 26314
rect 47952 26250 48004 26256
rect 47964 25945 47992 26250
rect 47950 25936 48006 25945
rect 47950 25871 48006 25880
rect 47872 25350 47992 25378
rect 47860 25288 47912 25294
rect 47858 25256 47860 25265
rect 47912 25256 47914 25265
rect 47858 25191 47914 25200
rect 47964 24018 47992 25350
rect 48056 24954 48084 27814
rect 48136 26308 48188 26314
rect 48136 26250 48188 26256
rect 48044 24948 48096 24954
rect 48044 24890 48096 24896
rect 48148 24682 48176 26250
rect 48136 24676 48188 24682
rect 48136 24618 48188 24624
rect 48134 24576 48190 24585
rect 48134 24511 48190 24520
rect 48044 24336 48096 24342
rect 48044 24278 48096 24284
rect 47872 23990 47992 24018
rect 47768 22228 47820 22234
rect 47768 22170 47820 22176
rect 47872 22114 47900 23990
rect 47950 23896 48006 23905
rect 48056 23866 48084 24278
rect 48148 24274 48176 24511
rect 48136 24268 48188 24274
rect 48136 24210 48188 24216
rect 47950 23831 48006 23840
rect 48044 23860 48096 23866
rect 47964 23798 47992 23831
rect 48044 23802 48096 23808
rect 47952 23792 48004 23798
rect 47952 23734 48004 23740
rect 48136 22636 48188 22642
rect 48136 22578 48188 22584
rect 48148 22545 48176 22578
rect 48134 22536 48190 22545
rect 48134 22471 48190 22480
rect 47780 22086 47900 22114
rect 47584 22024 47636 22030
rect 47584 21966 47636 21972
rect 47780 21690 47808 22086
rect 47860 22024 47912 22030
rect 47860 21966 47912 21972
rect 47768 21684 47820 21690
rect 47768 21626 47820 21632
rect 47768 19916 47820 19922
rect 47768 19858 47820 19864
rect 47780 19310 47808 19858
rect 47768 19304 47820 19310
rect 47768 19246 47820 19252
rect 47676 16992 47728 16998
rect 47676 16934 47728 16940
rect 47688 16522 47716 16934
rect 47676 16516 47728 16522
rect 47676 16458 47728 16464
rect 47872 15162 47900 21966
rect 47950 21856 48006 21865
rect 47950 21791 48006 21800
rect 47964 21622 47992 21791
rect 47952 21616 48004 21622
rect 47952 21558 48004 21564
rect 48044 21344 48096 21350
rect 48044 21286 48096 21292
rect 48056 20534 48084 21286
rect 48044 20528 48096 20534
rect 48044 20470 48096 20476
rect 48134 19816 48190 19825
rect 48134 19751 48136 19760
rect 48188 19751 48190 19760
rect 48136 19722 48188 19728
rect 48134 17096 48190 17105
rect 48134 17031 48190 17040
rect 48148 16658 48176 17031
rect 48136 16652 48188 16658
rect 48136 16594 48188 16600
rect 48134 16416 48190 16425
rect 48134 16351 48190 16360
rect 48148 15570 48176 16351
rect 48136 15564 48188 15570
rect 48136 15506 48188 15512
rect 47860 15156 47912 15162
rect 47860 15098 47912 15104
rect 47768 14816 47820 14822
rect 47768 14758 47820 14764
rect 47780 14482 47808 14758
rect 48044 14612 48096 14618
rect 48044 14554 48096 14560
rect 47768 14476 47820 14482
rect 47768 14418 47820 14424
rect 48056 14074 48084 14554
rect 48134 14376 48190 14385
rect 48134 14311 48136 14320
rect 48188 14311 48190 14320
rect 48136 14282 48188 14288
rect 48044 14068 48096 14074
rect 48044 14010 48096 14016
rect 47860 13932 47912 13938
rect 47860 13874 47912 13880
rect 47872 13705 47900 13874
rect 47858 13696 47914 13705
rect 47858 13631 47914 13640
rect 48136 11076 48188 11082
rect 48136 11018 48188 11024
rect 48148 10985 48176 11018
rect 48134 10976 48190 10985
rect 48134 10911 48190 10920
rect 47768 10668 47820 10674
rect 47768 10610 47820 10616
rect 47780 10305 47808 10610
rect 47766 10296 47822 10305
rect 47766 10231 47822 10240
rect 47950 8936 48006 8945
rect 47950 8871 47952 8880
rect 48004 8871 48006 8880
rect 47952 8842 48004 8848
rect 47768 8492 47820 8498
rect 47768 8434 47820 8440
rect 47780 8265 47808 8434
rect 47766 8256 47822 8265
rect 47766 8191 47822 8200
rect 48134 7576 48190 7585
rect 48134 7511 48190 7520
rect 47768 7200 47820 7206
rect 47768 7142 47820 7148
rect 47780 6730 47808 7142
rect 48148 6866 48176 7511
rect 48136 6860 48188 6866
rect 48136 6802 48188 6808
rect 47768 6724 47820 6730
rect 47768 6666 47820 6672
rect 47952 5636 48004 5642
rect 47952 5578 48004 5584
rect 47964 5545 47992 5578
rect 47950 5536 48006 5545
rect 47950 5471 48006 5480
rect 48240 5234 48268 35430
rect 48332 33318 48360 35550
rect 48320 33312 48372 33318
rect 48320 33254 48372 33260
rect 48504 30660 48556 30666
rect 48504 30602 48556 30608
rect 47492 5228 47544 5234
rect 47492 5170 47544 5176
rect 47584 5228 47636 5234
rect 47584 5170 47636 5176
rect 48228 5228 48280 5234
rect 48228 5170 48280 5176
rect 47400 4752 47452 4758
rect 47400 4694 47452 4700
rect 47596 3738 47624 5170
rect 47676 5024 47728 5030
rect 47676 4966 47728 4972
rect 47688 4690 47716 4966
rect 48134 4856 48190 4865
rect 48134 4791 48190 4800
rect 48148 4690 48176 4791
rect 47676 4684 47728 4690
rect 47676 4626 47728 4632
rect 48136 4684 48188 4690
rect 48136 4626 48188 4632
rect 48044 3936 48096 3942
rect 48044 3878 48096 3884
rect 47584 3732 47636 3738
rect 47584 3674 47636 3680
rect 47216 3460 47268 3466
rect 47216 3402 47268 3408
rect 48056 3194 48084 3878
rect 48044 3188 48096 3194
rect 48044 3130 48096 3136
rect 48320 2440 48372 2446
rect 48320 2382 48372 2388
rect 47768 2372 47820 2378
rect 47768 2314 47820 2320
rect 46754 96 46810 105
rect 46754 31 46810 40
rect 47030 0 47086 800
rect 47674 0 47730 800
rect 47780 785 47808 2314
rect 47860 2304 47912 2310
rect 47860 2246 47912 2252
rect 47872 1902 47900 2246
rect 47860 1896 47912 1902
rect 47860 1838 47912 1844
rect 48332 800 48360 2382
rect 47766 776 47822 785
rect 47766 711 47822 720
rect 48318 0 48374 800
rect 48516 762 48544 30602
rect 49608 3052 49660 3058
rect 49608 2994 49660 3000
rect 48884 870 49004 898
rect 48884 762 48912 870
rect 48976 800 49004 870
rect 49620 800 49648 2994
rect 48516 734 48912 762
rect 48962 0 49018 800
rect 49606 0 49662 800
<< via2 >>
rect 2870 51720 2926 51776
rect 1398 45600 1454 45656
rect 1398 40160 1454 40216
rect 1398 36760 1454 36816
rect 1398 34720 1454 34776
rect 1858 46960 1914 47016
rect 4066 51040 4122 51096
rect 3974 50360 4030 50416
rect 1490 31356 1492 31376
rect 1492 31356 1544 31376
rect 1544 31356 1546 31376
rect 1490 31320 1546 31356
rect 1398 23840 1454 23896
rect 1582 25900 1638 25936
rect 1582 25880 1584 25900
rect 1584 25880 1636 25900
rect 1636 25880 1638 25900
rect 2778 46280 2834 46336
rect 2778 44940 2834 44976
rect 2778 44920 2780 44940
rect 2780 44920 2832 44940
rect 2832 44920 2834 44940
rect 1858 44240 1914 44296
rect 1858 43560 1914 43616
rect 1858 41520 1914 41576
rect 1858 40840 1914 40896
rect 1858 37440 1914 37496
rect 3146 49000 3202 49056
rect 3422 48340 3478 48376
rect 3422 48320 3424 48340
rect 3424 48320 3476 48340
rect 3476 48320 3478 48340
rect 4220 49530 4276 49532
rect 4300 49530 4356 49532
rect 4380 49530 4436 49532
rect 4460 49530 4516 49532
rect 4220 49478 4266 49530
rect 4266 49478 4276 49530
rect 4300 49478 4330 49530
rect 4330 49478 4342 49530
rect 4342 49478 4356 49530
rect 4380 49478 4394 49530
rect 4394 49478 4406 49530
rect 4406 49478 4436 49530
rect 4460 49478 4470 49530
rect 4470 49478 4516 49530
rect 4220 49476 4276 49478
rect 4300 49476 4356 49478
rect 4380 49476 4436 49478
rect 4460 49476 4516 49478
rect 4220 48442 4276 48444
rect 4300 48442 4356 48444
rect 4380 48442 4436 48444
rect 4460 48442 4516 48444
rect 4220 48390 4266 48442
rect 4266 48390 4276 48442
rect 4300 48390 4330 48442
rect 4330 48390 4342 48442
rect 4342 48390 4356 48442
rect 4380 48390 4394 48442
rect 4394 48390 4406 48442
rect 4406 48390 4436 48442
rect 4460 48390 4470 48442
rect 4470 48390 4516 48442
rect 4220 48388 4276 48390
rect 4300 48388 4356 48390
rect 4380 48388 4436 48390
rect 4460 48388 4516 48390
rect 3790 47640 3846 47696
rect 2870 39480 2926 39536
rect 4220 47354 4276 47356
rect 4300 47354 4356 47356
rect 4380 47354 4436 47356
rect 4460 47354 4516 47356
rect 4220 47302 4266 47354
rect 4266 47302 4276 47354
rect 4300 47302 4330 47354
rect 4330 47302 4342 47354
rect 4342 47302 4356 47354
rect 4380 47302 4394 47354
rect 4394 47302 4406 47354
rect 4406 47302 4436 47354
rect 4460 47302 4470 47354
rect 4470 47302 4516 47354
rect 4220 47300 4276 47302
rect 4300 47300 4356 47302
rect 4380 47300 4436 47302
rect 4460 47300 4516 47302
rect 4220 46266 4276 46268
rect 4300 46266 4356 46268
rect 4380 46266 4436 46268
rect 4460 46266 4516 46268
rect 4220 46214 4266 46266
rect 4266 46214 4276 46266
rect 4300 46214 4330 46266
rect 4330 46214 4342 46266
rect 4342 46214 4356 46266
rect 4380 46214 4394 46266
rect 4394 46214 4406 46266
rect 4406 46214 4436 46266
rect 4460 46214 4470 46266
rect 4470 46214 4516 46266
rect 4220 46212 4276 46214
rect 4300 46212 4356 46214
rect 4380 46212 4436 46214
rect 4460 46212 4516 46214
rect 4220 45178 4276 45180
rect 4300 45178 4356 45180
rect 4380 45178 4436 45180
rect 4460 45178 4516 45180
rect 4220 45126 4266 45178
rect 4266 45126 4276 45178
rect 4300 45126 4330 45178
rect 4330 45126 4342 45178
rect 4342 45126 4356 45178
rect 4380 45126 4394 45178
rect 4394 45126 4406 45178
rect 4406 45126 4436 45178
rect 4460 45126 4470 45178
rect 4470 45126 4516 45178
rect 4220 45124 4276 45126
rect 4300 45124 4356 45126
rect 4380 45124 4436 45126
rect 4460 45124 4516 45126
rect 4220 44090 4276 44092
rect 4300 44090 4356 44092
rect 4380 44090 4436 44092
rect 4460 44090 4516 44092
rect 4220 44038 4266 44090
rect 4266 44038 4276 44090
rect 4300 44038 4330 44090
rect 4330 44038 4342 44090
rect 4342 44038 4356 44090
rect 4380 44038 4394 44090
rect 4394 44038 4406 44090
rect 4406 44038 4436 44090
rect 4460 44038 4470 44090
rect 4470 44038 4516 44090
rect 4220 44036 4276 44038
rect 4300 44036 4356 44038
rect 4380 44036 4436 44038
rect 4460 44036 4516 44038
rect 4220 43002 4276 43004
rect 4300 43002 4356 43004
rect 4380 43002 4436 43004
rect 4460 43002 4516 43004
rect 4220 42950 4266 43002
rect 4266 42950 4276 43002
rect 4300 42950 4330 43002
rect 4330 42950 4342 43002
rect 4342 42950 4356 43002
rect 4380 42950 4394 43002
rect 4394 42950 4406 43002
rect 4406 42950 4436 43002
rect 4460 42950 4470 43002
rect 4470 42950 4516 43002
rect 4220 42948 4276 42950
rect 4300 42948 4356 42950
rect 4380 42948 4436 42950
rect 4460 42948 4516 42950
rect 4220 41914 4276 41916
rect 4300 41914 4356 41916
rect 4380 41914 4436 41916
rect 4460 41914 4516 41916
rect 4220 41862 4266 41914
rect 4266 41862 4276 41914
rect 4300 41862 4330 41914
rect 4330 41862 4342 41914
rect 4342 41862 4356 41914
rect 4380 41862 4394 41914
rect 4394 41862 4406 41914
rect 4406 41862 4436 41914
rect 4460 41862 4470 41914
rect 4470 41862 4516 41914
rect 4220 41860 4276 41862
rect 4300 41860 4356 41862
rect 4380 41860 4436 41862
rect 4460 41860 4516 41862
rect 4220 40826 4276 40828
rect 4300 40826 4356 40828
rect 4380 40826 4436 40828
rect 4460 40826 4516 40828
rect 4220 40774 4266 40826
rect 4266 40774 4276 40826
rect 4300 40774 4330 40826
rect 4330 40774 4342 40826
rect 4342 40774 4356 40826
rect 4380 40774 4394 40826
rect 4394 40774 4406 40826
rect 4406 40774 4436 40826
rect 4460 40774 4470 40826
rect 4470 40774 4516 40826
rect 4220 40772 4276 40774
rect 4300 40772 4356 40774
rect 4380 40772 4436 40774
rect 4460 40772 4516 40774
rect 4220 39738 4276 39740
rect 4300 39738 4356 39740
rect 4380 39738 4436 39740
rect 4460 39738 4516 39740
rect 4220 39686 4266 39738
rect 4266 39686 4276 39738
rect 4300 39686 4330 39738
rect 4330 39686 4342 39738
rect 4342 39686 4356 39738
rect 4380 39686 4394 39738
rect 4394 39686 4406 39738
rect 4406 39686 4436 39738
rect 4460 39686 4470 39738
rect 4470 39686 4516 39738
rect 4220 39684 4276 39686
rect 4300 39684 4356 39686
rect 4380 39684 4436 39686
rect 4460 39684 4516 39686
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 4066 38120 4122 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 2778 36080 2834 36136
rect 1858 22480 1914 22536
rect 2778 34060 2834 34096
rect 2778 34040 2780 34060
rect 2780 34040 2832 34060
rect 2832 34040 2834 34060
rect 2778 33360 2834 33416
rect 1858 17040 1914 17096
rect 1398 12280 1454 12336
rect 1398 10920 1454 10976
rect 1858 8200 1914 8256
rect 1858 7520 1914 7576
rect 3146 32680 3202 32736
rect 3238 32000 3294 32056
rect 2778 29960 2834 30016
rect 2778 28620 2834 28656
rect 2778 28600 2780 28620
rect 2780 28600 2832 28620
rect 2832 28600 2834 28620
rect 2778 27240 2834 27296
rect 2778 26560 2834 26616
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4066 29280 4122 29336
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 1858 3440 1914 3496
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 2778 23180 2834 23216
rect 2778 23160 2780 23180
rect 2780 23160 2832 23180
rect 2832 23160 2834 23180
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 3974 21800 4030 21856
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4066 21120 4122 21176
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4066 19760 4122 19816
rect 2778 19080 2834 19136
rect 3146 18400 3202 18456
rect 2778 17740 2834 17776
rect 2778 17720 2780 17740
rect 2780 17720 2832 17740
rect 2832 17720 2834 17740
rect 2778 16360 2834 16416
rect 2778 13640 2834 13696
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 3054 10240 3110 10296
rect 3238 9560 3294 9616
rect 2962 8880 3018 8936
rect 2778 6860 2834 6896
rect 2778 6840 2780 6860
rect 2780 6840 2832 6860
rect 2832 6840 2834 6860
rect 3422 6160 3478 6216
rect 2778 5480 2834 5536
rect 3238 4800 3294 4856
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4066 12960 4122 13016
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 3422 4156 3424 4176
rect 3424 4156 3476 4176
rect 3476 4156 3478 4176
rect 3422 4120 3478 4156
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4066 2080 4122 2136
rect 4802 2352 4858 2408
rect 2778 720 2834 776
rect 11150 28736 11206 28792
rect 10322 23060 10324 23080
rect 10324 23060 10376 23080
rect 10376 23060 10378 23080
rect 10322 23024 10378 23060
rect 12070 28500 12072 28520
rect 12072 28500 12124 28520
rect 12124 28500 12126 28520
rect 12070 28464 12126 28500
rect 11978 23588 12034 23624
rect 11978 23568 11980 23588
rect 11980 23568 12032 23588
rect 12032 23568 12034 23588
rect 10966 20460 11022 20496
rect 10966 20440 10968 20460
rect 10968 20440 11020 20460
rect 11020 20440 11022 20460
rect 10966 18300 10968 18320
rect 10968 18300 11020 18320
rect 11020 18300 11022 18320
rect 10966 18264 11022 18300
rect 12990 31356 12992 31376
rect 12992 31356 13044 31376
rect 13044 31356 13046 31376
rect 12990 31320 13046 31356
rect 12714 25880 12770 25936
rect 14094 31320 14150 31376
rect 16670 47504 16726 47560
rect 17406 47524 17462 47560
rect 17406 47504 17408 47524
rect 17408 47504 17460 47524
rect 17460 47504 17462 47524
rect 19580 48986 19636 48988
rect 19660 48986 19716 48988
rect 19740 48986 19796 48988
rect 19820 48986 19876 48988
rect 19580 48934 19626 48986
rect 19626 48934 19636 48986
rect 19660 48934 19690 48986
rect 19690 48934 19702 48986
rect 19702 48934 19716 48986
rect 19740 48934 19754 48986
rect 19754 48934 19766 48986
rect 19766 48934 19796 48986
rect 19820 48934 19830 48986
rect 19830 48934 19876 48986
rect 19580 48932 19636 48934
rect 19660 48932 19716 48934
rect 19740 48932 19796 48934
rect 19820 48932 19876 48934
rect 13910 28600 13966 28656
rect 12438 20460 12494 20496
rect 12438 20440 12440 20460
rect 12440 20440 12492 20460
rect 12492 20440 12494 20460
rect 12254 20168 12310 20224
rect 11978 19896 12034 19952
rect 11978 19488 12034 19544
rect 12622 19760 12678 19816
rect 12254 18284 12310 18320
rect 12254 18264 12256 18284
rect 12256 18264 12308 18284
rect 12308 18264 12310 18284
rect 14278 25780 14280 25800
rect 14280 25780 14332 25800
rect 14332 25780 14334 25800
rect 14278 25744 14334 25780
rect 15658 28736 15714 28792
rect 16026 29008 16082 29064
rect 16762 28736 16818 28792
rect 15474 26308 15530 26344
rect 15474 26288 15476 26308
rect 15476 26288 15528 26308
rect 15528 26288 15530 26308
rect 16210 25608 16266 25664
rect 14462 23024 14518 23080
rect 13266 19488 13322 19544
rect 17682 28464 17738 28520
rect 19580 47898 19636 47900
rect 19660 47898 19716 47900
rect 19740 47898 19796 47900
rect 19820 47898 19876 47900
rect 19580 47846 19626 47898
rect 19626 47846 19636 47898
rect 19660 47846 19690 47898
rect 19690 47846 19702 47898
rect 19702 47846 19716 47898
rect 19740 47846 19754 47898
rect 19754 47846 19766 47898
rect 19766 47846 19796 47898
rect 19820 47846 19830 47898
rect 19830 47846 19876 47898
rect 19580 47844 19636 47846
rect 19660 47844 19716 47846
rect 19740 47844 19796 47846
rect 19820 47844 19876 47846
rect 19580 46810 19636 46812
rect 19660 46810 19716 46812
rect 19740 46810 19796 46812
rect 19820 46810 19876 46812
rect 19580 46758 19626 46810
rect 19626 46758 19636 46810
rect 19660 46758 19690 46810
rect 19690 46758 19702 46810
rect 19702 46758 19716 46810
rect 19740 46758 19754 46810
rect 19754 46758 19766 46810
rect 19766 46758 19796 46810
rect 19820 46758 19830 46810
rect 19830 46758 19876 46810
rect 19580 46756 19636 46758
rect 19660 46756 19716 46758
rect 19740 46756 19796 46758
rect 19820 46756 19876 46758
rect 19580 45722 19636 45724
rect 19660 45722 19716 45724
rect 19740 45722 19796 45724
rect 19820 45722 19876 45724
rect 19580 45670 19626 45722
rect 19626 45670 19636 45722
rect 19660 45670 19690 45722
rect 19690 45670 19702 45722
rect 19702 45670 19716 45722
rect 19740 45670 19754 45722
rect 19754 45670 19766 45722
rect 19766 45670 19796 45722
rect 19820 45670 19830 45722
rect 19830 45670 19876 45722
rect 19580 45668 19636 45670
rect 19660 45668 19716 45670
rect 19740 45668 19796 45670
rect 19820 45668 19876 45670
rect 19580 44634 19636 44636
rect 19660 44634 19716 44636
rect 19740 44634 19796 44636
rect 19820 44634 19876 44636
rect 19580 44582 19626 44634
rect 19626 44582 19636 44634
rect 19660 44582 19690 44634
rect 19690 44582 19702 44634
rect 19702 44582 19716 44634
rect 19740 44582 19754 44634
rect 19754 44582 19766 44634
rect 19766 44582 19796 44634
rect 19820 44582 19830 44634
rect 19830 44582 19876 44634
rect 19580 44580 19636 44582
rect 19660 44580 19716 44582
rect 19740 44580 19796 44582
rect 19820 44580 19876 44582
rect 19580 43546 19636 43548
rect 19660 43546 19716 43548
rect 19740 43546 19796 43548
rect 19820 43546 19876 43548
rect 19580 43494 19626 43546
rect 19626 43494 19636 43546
rect 19660 43494 19690 43546
rect 19690 43494 19702 43546
rect 19702 43494 19716 43546
rect 19740 43494 19754 43546
rect 19754 43494 19766 43546
rect 19766 43494 19796 43546
rect 19820 43494 19830 43546
rect 19830 43494 19876 43546
rect 19580 43492 19636 43494
rect 19660 43492 19716 43494
rect 19740 43492 19796 43494
rect 19820 43492 19876 43494
rect 19580 42458 19636 42460
rect 19660 42458 19716 42460
rect 19740 42458 19796 42460
rect 19820 42458 19876 42460
rect 19580 42406 19626 42458
rect 19626 42406 19636 42458
rect 19660 42406 19690 42458
rect 19690 42406 19702 42458
rect 19702 42406 19716 42458
rect 19740 42406 19754 42458
rect 19754 42406 19766 42458
rect 19766 42406 19796 42458
rect 19820 42406 19830 42458
rect 19830 42406 19876 42458
rect 19580 42404 19636 42406
rect 19660 42404 19716 42406
rect 19740 42404 19796 42406
rect 19820 42404 19876 42406
rect 19580 41370 19636 41372
rect 19660 41370 19716 41372
rect 19740 41370 19796 41372
rect 19820 41370 19876 41372
rect 19580 41318 19626 41370
rect 19626 41318 19636 41370
rect 19660 41318 19690 41370
rect 19690 41318 19702 41370
rect 19702 41318 19716 41370
rect 19740 41318 19754 41370
rect 19754 41318 19766 41370
rect 19766 41318 19796 41370
rect 19820 41318 19830 41370
rect 19830 41318 19876 41370
rect 19580 41316 19636 41318
rect 19660 41316 19716 41318
rect 19740 41316 19796 41318
rect 19820 41316 19876 41318
rect 19580 40282 19636 40284
rect 19660 40282 19716 40284
rect 19740 40282 19796 40284
rect 19820 40282 19876 40284
rect 19580 40230 19626 40282
rect 19626 40230 19636 40282
rect 19660 40230 19690 40282
rect 19690 40230 19702 40282
rect 19702 40230 19716 40282
rect 19740 40230 19754 40282
rect 19754 40230 19766 40282
rect 19766 40230 19796 40282
rect 19820 40230 19830 40282
rect 19830 40230 19876 40282
rect 19580 40228 19636 40230
rect 19660 40228 19716 40230
rect 19740 40228 19796 40230
rect 19820 40228 19876 40230
rect 19580 39194 19636 39196
rect 19660 39194 19716 39196
rect 19740 39194 19796 39196
rect 19820 39194 19876 39196
rect 19580 39142 19626 39194
rect 19626 39142 19636 39194
rect 19660 39142 19690 39194
rect 19690 39142 19702 39194
rect 19702 39142 19716 39194
rect 19740 39142 19754 39194
rect 19754 39142 19766 39194
rect 19766 39142 19796 39194
rect 19820 39142 19830 39194
rect 19830 39142 19876 39194
rect 19580 39140 19636 39142
rect 19660 39140 19716 39142
rect 19740 39140 19796 39142
rect 19820 39140 19876 39142
rect 18050 29028 18106 29064
rect 18050 29008 18052 29028
rect 18052 29008 18104 29028
rect 18104 29008 18106 29028
rect 18142 28600 18198 28656
rect 17682 26288 17738 26344
rect 17130 25744 17186 25800
rect 17406 25916 17408 25936
rect 17408 25916 17460 25936
rect 17460 25916 17462 25936
rect 17406 25880 17462 25916
rect 18234 25644 18236 25664
rect 18236 25644 18288 25664
rect 18288 25644 18290 25664
rect 14278 19896 14334 19952
rect 15934 20340 15936 20360
rect 15936 20340 15988 20360
rect 15988 20340 15990 20360
rect 15934 20304 15990 20340
rect 12438 4020 12440 4040
rect 12440 4020 12492 4040
rect 12492 4020 12494 4040
rect 12438 3984 12494 4020
rect 18234 25608 18290 25644
rect 18050 23724 18106 23760
rect 18050 23704 18052 23724
rect 18052 23704 18104 23724
rect 18104 23704 18106 23724
rect 18418 23604 18420 23624
rect 18420 23604 18472 23624
rect 18472 23604 18474 23624
rect 18418 23568 18474 23604
rect 17682 22480 17738 22536
rect 17498 20168 17554 20224
rect 17682 19796 17684 19816
rect 17684 19796 17736 19816
rect 17736 19796 17738 19816
rect 17682 19760 17738 19796
rect 18234 19488 18290 19544
rect 18602 20304 18658 20360
rect 18694 19796 18696 19816
rect 18696 19796 18748 19816
rect 18748 19796 18750 19816
rect 18694 19760 18750 19796
rect 17682 3984 17738 4040
rect 19580 38106 19636 38108
rect 19660 38106 19716 38108
rect 19740 38106 19796 38108
rect 19820 38106 19876 38108
rect 19580 38054 19626 38106
rect 19626 38054 19636 38106
rect 19660 38054 19690 38106
rect 19690 38054 19702 38106
rect 19702 38054 19716 38106
rect 19740 38054 19754 38106
rect 19754 38054 19766 38106
rect 19766 38054 19796 38106
rect 19820 38054 19830 38106
rect 19830 38054 19876 38106
rect 19580 38052 19636 38054
rect 19660 38052 19716 38054
rect 19740 38052 19796 38054
rect 19820 38052 19876 38054
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19798 35436 19800 35456
rect 19800 35436 19852 35456
rect 19852 35436 19854 35456
rect 19798 35400 19854 35436
rect 19614 35128 19670 35184
rect 19890 34992 19946 35048
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19522 29144 19578 29200
rect 20258 40704 20314 40760
rect 20166 32952 20222 33008
rect 20350 40432 20406 40488
rect 20258 30776 20314 30832
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19706 27412 19708 27432
rect 19708 27412 19760 27432
rect 19760 27412 19762 27432
rect 19706 27376 19762 27412
rect 20074 27376 20130 27432
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 20074 24928 20130 24984
rect 19982 24656 20038 24712
rect 19890 24248 19946 24304
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19062 19488 19118 19544
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 20074 24384 20130 24440
rect 20442 38800 20498 38856
rect 20350 24792 20406 24848
rect 20350 24520 20406 24576
rect 20350 23604 20352 23624
rect 20352 23604 20404 23624
rect 20404 23604 20406 23624
rect 20350 23568 20406 23604
rect 20258 21956 20314 21992
rect 20258 21936 20260 21956
rect 20260 21936 20312 21956
rect 20312 21936 20314 21956
rect 20166 17448 20222 17504
rect 20350 17312 20406 17368
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 20718 39380 20720 39400
rect 20720 39380 20772 39400
rect 20772 39380 20774 39400
rect 20718 39344 20774 39380
rect 20902 38800 20958 38856
rect 20718 35708 20720 35728
rect 20720 35708 20772 35728
rect 20772 35708 20774 35728
rect 20718 35672 20774 35708
rect 20810 28364 20812 28384
rect 20812 28364 20864 28384
rect 20864 28364 20866 28384
rect 20810 28328 20866 28364
rect 20718 21528 20774 21584
rect 20626 18284 20682 18320
rect 20626 18264 20628 18284
rect 20628 18264 20680 18284
rect 20680 18264 20682 18284
rect 22282 38836 22284 38856
rect 22284 38836 22336 38856
rect 22336 38836 22338 38856
rect 22282 38800 22338 38836
rect 22374 36080 22430 36136
rect 21914 35692 21970 35728
rect 21914 35672 21916 35692
rect 21916 35672 21968 35692
rect 21968 35672 21970 35692
rect 22006 35400 22062 35456
rect 21454 34992 21510 35048
rect 21914 35028 21916 35048
rect 21916 35028 21968 35048
rect 21968 35028 21970 35048
rect 21914 34992 21970 35028
rect 21086 30232 21142 30288
rect 20994 21664 21050 21720
rect 21178 24384 21234 24440
rect 21178 21528 21234 21584
rect 21362 24656 21418 24712
rect 21638 24520 21694 24576
rect 22374 33496 22430 33552
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 21822 17856 21878 17912
rect 22098 21936 22154 21992
rect 23110 25064 23166 25120
rect 22926 24556 22928 24576
rect 22928 24556 22980 24576
rect 22980 24556 22982 24576
rect 22926 24520 22982 24556
rect 22098 18420 22154 18456
rect 22098 18400 22100 18420
rect 22100 18400 22152 18420
rect 22152 18400 22154 18420
rect 22466 17060 22522 17096
rect 22466 17040 22468 17060
rect 22468 17040 22520 17060
rect 22520 17040 22522 17060
rect 22374 16632 22430 16688
rect 22650 17448 22706 17504
rect 22558 3984 22614 4040
rect 22926 17312 22982 17368
rect 22926 16088 22982 16144
rect 23386 26968 23442 27024
rect 23754 27240 23810 27296
rect 24582 35128 24638 35184
rect 24030 33516 24086 33552
rect 24030 33496 24032 33516
rect 24032 33496 24084 33516
rect 24084 33496 24086 33516
rect 23846 24112 23902 24168
rect 23570 22480 23626 22536
rect 23294 20460 23350 20496
rect 23294 20440 23296 20460
rect 23296 20440 23348 20460
rect 23348 20440 23350 20460
rect 23202 20304 23258 20360
rect 23386 17584 23442 17640
rect 23386 17448 23442 17504
rect 23386 16768 23442 16824
rect 23478 16516 23534 16552
rect 23478 16496 23480 16516
rect 23480 16496 23532 16516
rect 23532 16496 23534 16516
rect 24490 25064 24546 25120
rect 25410 33516 25466 33552
rect 25410 33496 25412 33516
rect 25412 33496 25464 33516
rect 25464 33496 25466 33516
rect 26238 35572 26240 35592
rect 26240 35572 26292 35592
rect 26292 35572 26294 35592
rect 26238 35536 26294 35572
rect 25778 30776 25834 30832
rect 24674 24928 24730 24984
rect 24214 24520 24270 24576
rect 24674 24148 24676 24168
rect 24676 24148 24728 24168
rect 24728 24148 24730 24168
rect 24674 24112 24730 24148
rect 24582 23976 24638 24032
rect 23662 17060 23718 17096
rect 23662 17040 23664 17060
rect 23664 17040 23716 17060
rect 23716 17040 23718 17060
rect 23662 16108 23718 16144
rect 23662 16088 23664 16108
rect 23664 16088 23716 16108
rect 23716 16088 23718 16108
rect 23846 16632 23902 16688
rect 24398 22888 24454 22944
rect 24582 21836 24584 21856
rect 24584 21836 24636 21856
rect 24636 21836 24638 21856
rect 24582 21800 24638 21836
rect 24582 21664 24638 21720
rect 24398 20712 24454 20768
rect 25870 24556 25872 24576
rect 25872 24556 25924 24576
rect 25924 24556 25926 24576
rect 25870 24520 25926 24556
rect 25686 19352 25742 19408
rect 25318 18284 25374 18320
rect 25318 18264 25320 18284
rect 25320 18264 25372 18284
rect 25372 18264 25374 18284
rect 25686 18128 25742 18184
rect 26238 23568 26294 23624
rect 26238 20440 26294 20496
rect 26330 19216 26386 19272
rect 26054 18264 26110 18320
rect 26146 16088 26202 16144
rect 26606 39344 26662 39400
rect 26606 24248 26662 24304
rect 26238 12688 26294 12744
rect 24398 4004 24454 4040
rect 24398 3984 24400 4004
rect 24400 3984 24452 4004
rect 24452 3984 24454 4004
rect 27526 36116 27528 36136
rect 27528 36116 27580 36136
rect 27580 36116 27582 36136
rect 27526 36080 27582 36116
rect 27618 35536 27674 35592
rect 27158 33532 27160 33552
rect 27160 33532 27212 33552
rect 27212 33532 27214 33552
rect 27158 33496 27214 33532
rect 27434 28076 27490 28112
rect 27434 28056 27436 28076
rect 27436 28056 27488 28076
rect 27488 28056 27490 28076
rect 27434 26988 27490 27024
rect 27434 26968 27436 26988
rect 27436 26968 27488 26988
rect 27488 26968 27490 26988
rect 27158 24928 27214 24984
rect 27250 12688 27306 12744
rect 26790 9968 26846 10024
rect 27894 28328 27950 28384
rect 28078 28056 28134 28112
rect 27986 27240 28042 27296
rect 27802 21800 27858 21856
rect 27618 15680 27674 15736
rect 27802 15680 27858 15736
rect 28170 18400 28226 18456
rect 28170 17720 28226 17776
rect 28446 17856 28502 17912
rect 28354 16360 28410 16416
rect 28630 27276 28632 27296
rect 28632 27276 28684 27296
rect 28684 27276 28686 27296
rect 28630 27240 28686 27276
rect 29274 30232 29330 30288
rect 29274 28076 29330 28112
rect 29274 28056 29276 28076
rect 29276 28056 29328 28076
rect 29328 28056 29330 28076
rect 29550 26696 29606 26752
rect 28906 23976 28962 24032
rect 29550 15816 29606 15872
rect 28998 11056 29054 11112
rect 28998 10376 29054 10432
rect 28906 10004 28908 10024
rect 28908 10004 28960 10024
rect 28960 10004 28962 10024
rect 28906 9968 28962 10004
rect 29366 10412 29368 10432
rect 29368 10412 29420 10432
rect 29420 10412 29422 10432
rect 29366 10376 29422 10412
rect 30010 15952 30066 16008
rect 30286 15952 30342 16008
rect 30746 15680 30802 15736
rect 31022 15988 31024 16008
rect 31024 15988 31076 16008
rect 31076 15988 31078 16008
rect 31022 15952 31078 15988
rect 32402 26696 32458 26752
rect 33230 30252 33286 30288
rect 33230 30232 33232 30252
rect 33232 30232 33284 30252
rect 33284 30232 33286 30252
rect 32310 15852 32312 15872
rect 32312 15852 32364 15872
rect 32364 15852 32366 15872
rect 32310 15816 32366 15852
rect 30930 10376 30986 10432
rect 30194 2896 30250 2952
rect 31298 2932 31300 2952
rect 31300 2932 31352 2952
rect 31352 2932 31354 2952
rect 31298 2896 31354 2932
rect 34940 49530 34996 49532
rect 35020 49530 35076 49532
rect 35100 49530 35156 49532
rect 35180 49530 35236 49532
rect 34940 49478 34986 49530
rect 34986 49478 34996 49530
rect 35020 49478 35050 49530
rect 35050 49478 35062 49530
rect 35062 49478 35076 49530
rect 35100 49478 35114 49530
rect 35114 49478 35126 49530
rect 35126 49478 35156 49530
rect 35180 49478 35190 49530
rect 35190 49478 35236 49530
rect 34940 49476 34996 49478
rect 35020 49476 35076 49478
rect 35100 49476 35156 49478
rect 35180 49476 35236 49478
rect 34940 48442 34996 48444
rect 35020 48442 35076 48444
rect 35100 48442 35156 48444
rect 35180 48442 35236 48444
rect 34940 48390 34986 48442
rect 34986 48390 34996 48442
rect 35020 48390 35050 48442
rect 35050 48390 35062 48442
rect 35062 48390 35076 48442
rect 35100 48390 35114 48442
rect 35114 48390 35126 48442
rect 35126 48390 35156 48442
rect 35180 48390 35190 48442
rect 35190 48390 35236 48442
rect 34940 48388 34996 48390
rect 35020 48388 35076 48390
rect 35100 48388 35156 48390
rect 35180 48388 35236 48390
rect 34940 47354 34996 47356
rect 35020 47354 35076 47356
rect 35100 47354 35156 47356
rect 35180 47354 35236 47356
rect 34940 47302 34986 47354
rect 34986 47302 34996 47354
rect 35020 47302 35050 47354
rect 35050 47302 35062 47354
rect 35062 47302 35076 47354
rect 35100 47302 35114 47354
rect 35114 47302 35126 47354
rect 35126 47302 35156 47354
rect 35180 47302 35190 47354
rect 35190 47302 35236 47354
rect 34940 47300 34996 47302
rect 35020 47300 35076 47302
rect 35100 47300 35156 47302
rect 35180 47300 35236 47302
rect 34940 46266 34996 46268
rect 35020 46266 35076 46268
rect 35100 46266 35156 46268
rect 35180 46266 35236 46268
rect 34940 46214 34986 46266
rect 34986 46214 34996 46266
rect 35020 46214 35050 46266
rect 35050 46214 35062 46266
rect 35062 46214 35076 46266
rect 35100 46214 35114 46266
rect 35114 46214 35126 46266
rect 35126 46214 35156 46266
rect 35180 46214 35190 46266
rect 35190 46214 35236 46266
rect 34940 46212 34996 46214
rect 35020 46212 35076 46214
rect 35100 46212 35156 46214
rect 35180 46212 35236 46214
rect 34940 45178 34996 45180
rect 35020 45178 35076 45180
rect 35100 45178 35156 45180
rect 35180 45178 35236 45180
rect 34940 45126 34986 45178
rect 34986 45126 34996 45178
rect 35020 45126 35050 45178
rect 35050 45126 35062 45178
rect 35062 45126 35076 45178
rect 35100 45126 35114 45178
rect 35114 45126 35126 45178
rect 35126 45126 35156 45178
rect 35180 45126 35190 45178
rect 35190 45126 35236 45178
rect 34940 45124 34996 45126
rect 35020 45124 35076 45126
rect 35100 45124 35156 45126
rect 35180 45124 35236 45126
rect 34940 44090 34996 44092
rect 35020 44090 35076 44092
rect 35100 44090 35156 44092
rect 35180 44090 35236 44092
rect 34940 44038 34986 44090
rect 34986 44038 34996 44090
rect 35020 44038 35050 44090
rect 35050 44038 35062 44090
rect 35062 44038 35076 44090
rect 35100 44038 35114 44090
rect 35114 44038 35126 44090
rect 35126 44038 35156 44090
rect 35180 44038 35190 44090
rect 35190 44038 35236 44090
rect 34940 44036 34996 44038
rect 35020 44036 35076 44038
rect 35100 44036 35156 44038
rect 35180 44036 35236 44038
rect 34940 43002 34996 43004
rect 35020 43002 35076 43004
rect 35100 43002 35156 43004
rect 35180 43002 35236 43004
rect 34940 42950 34986 43002
rect 34986 42950 34996 43002
rect 35020 42950 35050 43002
rect 35050 42950 35062 43002
rect 35062 42950 35076 43002
rect 35100 42950 35114 43002
rect 35114 42950 35126 43002
rect 35126 42950 35156 43002
rect 35180 42950 35190 43002
rect 35190 42950 35236 43002
rect 34940 42948 34996 42950
rect 35020 42948 35076 42950
rect 35100 42948 35156 42950
rect 35180 42948 35236 42950
rect 34940 41914 34996 41916
rect 35020 41914 35076 41916
rect 35100 41914 35156 41916
rect 35180 41914 35236 41916
rect 34940 41862 34986 41914
rect 34986 41862 34996 41914
rect 35020 41862 35050 41914
rect 35050 41862 35062 41914
rect 35062 41862 35076 41914
rect 35100 41862 35114 41914
rect 35114 41862 35126 41914
rect 35126 41862 35156 41914
rect 35180 41862 35190 41914
rect 35190 41862 35236 41914
rect 34940 41860 34996 41862
rect 35020 41860 35076 41862
rect 35100 41860 35156 41862
rect 35180 41860 35236 41862
rect 34940 40826 34996 40828
rect 35020 40826 35076 40828
rect 35100 40826 35156 40828
rect 35180 40826 35236 40828
rect 34940 40774 34986 40826
rect 34986 40774 34996 40826
rect 35020 40774 35050 40826
rect 35050 40774 35062 40826
rect 35062 40774 35076 40826
rect 35100 40774 35114 40826
rect 35114 40774 35126 40826
rect 35126 40774 35156 40826
rect 35180 40774 35190 40826
rect 35190 40774 35236 40826
rect 34940 40772 34996 40774
rect 35020 40772 35076 40774
rect 35100 40772 35156 40774
rect 35180 40772 35236 40774
rect 34940 39738 34996 39740
rect 35020 39738 35076 39740
rect 35100 39738 35156 39740
rect 35180 39738 35236 39740
rect 34940 39686 34986 39738
rect 34986 39686 34996 39738
rect 35020 39686 35050 39738
rect 35050 39686 35062 39738
rect 35062 39686 35076 39738
rect 35100 39686 35114 39738
rect 35114 39686 35126 39738
rect 35126 39686 35156 39738
rect 35180 39686 35190 39738
rect 35190 39686 35236 39738
rect 34940 39684 34996 39686
rect 35020 39684 35076 39686
rect 35100 39684 35156 39686
rect 35180 39684 35236 39686
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 38106 24792 38162 24848
rect 35070 2524 35072 2544
rect 35072 2524 35124 2544
rect 35124 2524 35126 2544
rect 35070 2488 35126 2524
rect 46570 51720 46626 51776
rect 45558 51040 45614 51096
rect 45558 44920 45614 44976
rect 46846 50360 46902 50416
rect 46754 49680 46810 49736
rect 45558 26560 45614 26616
rect 46018 44260 46074 44296
rect 46018 44240 46020 44260
rect 46020 44240 46072 44260
rect 46072 44240 46074 44260
rect 46846 46960 46902 47016
rect 46846 37440 46902 37496
rect 46846 29280 46902 29336
rect 47766 49000 47822 49056
rect 47766 48320 47822 48376
rect 47306 40840 47362 40896
rect 47306 29960 47362 30016
rect 45650 17720 45706 17776
rect 44822 16768 44878 16824
rect 45650 16768 45706 16824
rect 45558 12280 45614 12336
rect 45558 6840 45614 6896
rect 45650 6160 45706 6216
rect 45558 3440 45614 3496
rect 47490 32000 47546 32056
rect 47306 19080 47362 19136
rect 46846 15020 46902 15056
rect 46846 15000 46848 15020
rect 46848 15000 46900 15020
rect 46900 15000 46902 15020
rect 46846 12960 46902 13016
rect 46386 9560 46442 9616
rect 46202 4120 46258 4176
rect 46846 1400 46902 1456
rect 47582 23704 47638 23760
rect 48134 46280 48190 46336
rect 48134 45600 48190 45656
rect 48134 43560 48190 43616
rect 47858 42880 47914 42936
rect 47950 42200 48006 42256
rect 48134 41540 48190 41576
rect 48134 41520 48136 41540
rect 48136 41520 48188 41540
rect 48188 41520 48190 41540
rect 48134 40160 48190 40216
rect 48226 39480 48282 39536
rect 47950 38800 48006 38856
rect 47858 38120 47914 38176
rect 47858 36116 47860 36136
rect 47860 36116 47912 36136
rect 47912 36116 47914 36136
rect 47858 36080 47914 36116
rect 48134 36760 48190 36816
rect 48134 35400 48190 35456
rect 48134 34720 48190 34776
rect 48042 34040 48098 34096
rect 47950 33360 48006 33416
rect 47950 31340 48006 31376
rect 47950 31320 47952 31340
rect 47952 31320 48004 31340
rect 48004 31320 48006 31340
rect 47858 27920 47914 27976
rect 48134 28620 48190 28656
rect 48134 28600 48136 28620
rect 48136 28600 48188 28620
rect 48188 28600 48190 28620
rect 47950 25880 48006 25936
rect 47858 25236 47860 25256
rect 47860 25236 47912 25256
rect 47912 25236 47914 25256
rect 47858 25200 47914 25236
rect 48134 24520 48190 24576
rect 47950 23840 48006 23896
rect 48134 22480 48190 22536
rect 47950 21800 48006 21856
rect 48134 19780 48190 19816
rect 48134 19760 48136 19780
rect 48136 19760 48188 19780
rect 48188 19760 48190 19780
rect 48134 17040 48190 17096
rect 48134 16360 48190 16416
rect 48134 14340 48190 14376
rect 48134 14320 48136 14340
rect 48136 14320 48188 14340
rect 48188 14320 48190 14340
rect 47858 13640 47914 13696
rect 48134 10920 48190 10976
rect 47766 10240 47822 10296
rect 47950 8900 48006 8936
rect 47950 8880 47952 8900
rect 47952 8880 48004 8900
rect 48004 8880 48006 8900
rect 47766 8200 47822 8256
rect 48134 7520 48190 7576
rect 47950 5480 48006 5536
rect 48134 4800 48190 4856
rect 46754 40 46810 96
rect 47766 720 47822 776
<< metal3 >>
rect 0 51778 800 51808
rect 2865 51778 2931 51781
rect 0 51776 2931 51778
rect 0 51720 2870 51776
rect 2926 51720 2931 51776
rect 0 51718 2931 51720
rect 0 51688 800 51718
rect 2865 51715 2931 51718
rect 46565 51778 46631 51781
rect 49200 51778 50000 51808
rect 46565 51776 50000 51778
rect 46565 51720 46570 51776
rect 46626 51720 50000 51776
rect 46565 51718 50000 51720
rect 46565 51715 46631 51718
rect 49200 51688 50000 51718
rect 0 51098 800 51128
rect 4061 51098 4127 51101
rect 0 51096 4127 51098
rect 0 51040 4066 51096
rect 4122 51040 4127 51096
rect 0 51038 4127 51040
rect 0 51008 800 51038
rect 4061 51035 4127 51038
rect 45553 51098 45619 51101
rect 49200 51098 50000 51128
rect 45553 51096 50000 51098
rect 45553 51040 45558 51096
rect 45614 51040 50000 51096
rect 45553 51038 50000 51040
rect 45553 51035 45619 51038
rect 49200 51008 50000 51038
rect 0 50418 800 50448
rect 3969 50418 4035 50421
rect 0 50416 4035 50418
rect 0 50360 3974 50416
rect 4030 50360 4035 50416
rect 0 50358 4035 50360
rect 0 50328 800 50358
rect 3969 50355 4035 50358
rect 46841 50418 46907 50421
rect 49200 50418 50000 50448
rect 46841 50416 50000 50418
rect 46841 50360 46846 50416
rect 46902 50360 50000 50416
rect 46841 50358 50000 50360
rect 46841 50355 46907 50358
rect 49200 50328 50000 50358
rect 0 49648 800 49768
rect 46749 49738 46815 49741
rect 49200 49738 50000 49768
rect 46749 49736 50000 49738
rect 46749 49680 46754 49736
rect 46810 49680 50000 49736
rect 46749 49678 50000 49680
rect 46749 49675 46815 49678
rect 49200 49648 50000 49678
rect 4208 49536 4528 49537
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 49471 4528 49472
rect 34928 49536 35248 49537
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 49471 35248 49472
rect 0 49058 800 49088
rect 3141 49058 3207 49061
rect 0 49056 3207 49058
rect 0 49000 3146 49056
rect 3202 49000 3207 49056
rect 0 48998 3207 49000
rect 0 48968 800 48998
rect 3141 48995 3207 48998
rect 47761 49058 47827 49061
rect 49200 49058 50000 49088
rect 47761 49056 50000 49058
rect 47761 49000 47766 49056
rect 47822 49000 50000 49056
rect 47761 48998 50000 49000
rect 47761 48995 47827 48998
rect 19568 48992 19888 48993
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 49200 48968 50000 48998
rect 19568 48927 19888 48928
rect 4208 48448 4528 48449
rect 0 48378 800 48408
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 48383 4528 48384
rect 34928 48448 35248 48449
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 48383 35248 48384
rect 3417 48378 3483 48381
rect 0 48376 3483 48378
rect 0 48320 3422 48376
rect 3478 48320 3483 48376
rect 0 48318 3483 48320
rect 0 48288 800 48318
rect 3417 48315 3483 48318
rect 47761 48378 47827 48381
rect 49200 48378 50000 48408
rect 47761 48376 50000 48378
rect 47761 48320 47766 48376
rect 47822 48320 50000 48376
rect 47761 48318 50000 48320
rect 47761 48315 47827 48318
rect 49200 48288 50000 48318
rect 19568 47904 19888 47905
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 47839 19888 47840
rect 0 47698 800 47728
rect 3785 47698 3851 47701
rect 0 47696 3851 47698
rect 0 47640 3790 47696
rect 3846 47640 3851 47696
rect 0 47638 3851 47640
rect 0 47608 800 47638
rect 3785 47635 3851 47638
rect 49200 47608 50000 47728
rect 16665 47562 16731 47565
rect 17401 47562 17467 47565
rect 16665 47560 17467 47562
rect 16665 47504 16670 47560
rect 16726 47504 17406 47560
rect 17462 47504 17467 47560
rect 16665 47502 17467 47504
rect 16665 47499 16731 47502
rect 17401 47499 17467 47502
rect 4208 47360 4528 47361
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 47295 4528 47296
rect 34928 47360 35248 47361
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 47295 35248 47296
rect 0 47018 800 47048
rect 1853 47018 1919 47021
rect 0 47016 1919 47018
rect 0 46960 1858 47016
rect 1914 46960 1919 47016
rect 0 46958 1919 46960
rect 0 46928 800 46958
rect 1853 46955 1919 46958
rect 46841 47018 46907 47021
rect 49200 47018 50000 47048
rect 46841 47016 50000 47018
rect 46841 46960 46846 47016
rect 46902 46960 50000 47016
rect 46841 46958 50000 46960
rect 46841 46955 46907 46958
rect 49200 46928 50000 46958
rect 19568 46816 19888 46817
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 46751 19888 46752
rect 0 46338 800 46368
rect 2773 46338 2839 46341
rect 0 46336 2839 46338
rect 0 46280 2778 46336
rect 2834 46280 2839 46336
rect 0 46278 2839 46280
rect 0 46248 800 46278
rect 2773 46275 2839 46278
rect 48129 46338 48195 46341
rect 49200 46338 50000 46368
rect 48129 46336 50000 46338
rect 48129 46280 48134 46336
rect 48190 46280 50000 46336
rect 48129 46278 50000 46280
rect 48129 46275 48195 46278
rect 4208 46272 4528 46273
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 46207 4528 46208
rect 34928 46272 35248 46273
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 49200 46248 50000 46278
rect 34928 46207 35248 46208
rect 19568 45728 19888 45729
rect 0 45658 800 45688
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 45663 19888 45664
rect 1393 45658 1459 45661
rect 0 45656 1459 45658
rect 0 45600 1398 45656
rect 1454 45600 1459 45656
rect 0 45598 1459 45600
rect 0 45568 800 45598
rect 1393 45595 1459 45598
rect 48129 45658 48195 45661
rect 49200 45658 50000 45688
rect 48129 45656 50000 45658
rect 48129 45600 48134 45656
rect 48190 45600 50000 45656
rect 48129 45598 50000 45600
rect 48129 45595 48195 45598
rect 49200 45568 50000 45598
rect 4208 45184 4528 45185
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 45119 4528 45120
rect 34928 45184 35248 45185
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 45119 35248 45120
rect 0 44978 800 45008
rect 2773 44978 2839 44981
rect 0 44976 2839 44978
rect 0 44920 2778 44976
rect 2834 44920 2839 44976
rect 0 44918 2839 44920
rect 0 44888 800 44918
rect 2773 44915 2839 44918
rect 45553 44978 45619 44981
rect 49200 44978 50000 45008
rect 45553 44976 50000 44978
rect 45553 44920 45558 44976
rect 45614 44920 50000 44976
rect 45553 44918 50000 44920
rect 45553 44915 45619 44918
rect 49200 44888 50000 44918
rect 19568 44640 19888 44641
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 44575 19888 44576
rect 0 44298 800 44328
rect 1853 44298 1919 44301
rect 0 44296 1919 44298
rect 0 44240 1858 44296
rect 1914 44240 1919 44296
rect 0 44238 1919 44240
rect 0 44208 800 44238
rect 1853 44235 1919 44238
rect 46013 44298 46079 44301
rect 49200 44298 50000 44328
rect 46013 44296 50000 44298
rect 46013 44240 46018 44296
rect 46074 44240 50000 44296
rect 46013 44238 50000 44240
rect 46013 44235 46079 44238
rect 49200 44208 50000 44238
rect 4208 44096 4528 44097
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 44031 4528 44032
rect 34928 44096 35248 44097
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 44031 35248 44032
rect 0 43618 800 43648
rect 1853 43618 1919 43621
rect 0 43616 1919 43618
rect 0 43560 1858 43616
rect 1914 43560 1919 43616
rect 0 43558 1919 43560
rect 0 43528 800 43558
rect 1853 43555 1919 43558
rect 48129 43618 48195 43621
rect 49200 43618 50000 43648
rect 48129 43616 50000 43618
rect 48129 43560 48134 43616
rect 48190 43560 50000 43616
rect 48129 43558 50000 43560
rect 48129 43555 48195 43558
rect 19568 43552 19888 43553
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 49200 43528 50000 43558
rect 19568 43487 19888 43488
rect 4208 43008 4528 43009
rect 0 42848 800 42968
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 42943 4528 42944
rect 34928 43008 35248 43009
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 42943 35248 42944
rect 47853 42938 47919 42941
rect 49200 42938 50000 42968
rect 47853 42936 50000 42938
rect 47853 42880 47858 42936
rect 47914 42880 50000 42936
rect 47853 42878 50000 42880
rect 47853 42875 47919 42878
rect 49200 42848 50000 42878
rect 19568 42464 19888 42465
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 42399 19888 42400
rect 47945 42258 48011 42261
rect 49200 42258 50000 42288
rect 47945 42256 50000 42258
rect 47945 42200 47950 42256
rect 48006 42200 50000 42256
rect 47945 42198 50000 42200
rect 47945 42195 48011 42198
rect 49200 42168 50000 42198
rect 4208 41920 4528 41921
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 41855 4528 41856
rect 34928 41920 35248 41921
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 41855 35248 41856
rect 0 41578 800 41608
rect 1853 41578 1919 41581
rect 0 41576 1919 41578
rect 0 41520 1858 41576
rect 1914 41520 1919 41576
rect 0 41518 1919 41520
rect 0 41488 800 41518
rect 1853 41515 1919 41518
rect 48129 41578 48195 41581
rect 49200 41578 50000 41608
rect 48129 41576 50000 41578
rect 48129 41520 48134 41576
rect 48190 41520 50000 41576
rect 48129 41518 50000 41520
rect 48129 41515 48195 41518
rect 49200 41488 50000 41518
rect 19568 41376 19888 41377
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 41311 19888 41312
rect 0 40898 800 40928
rect 1853 40898 1919 40901
rect 0 40896 1919 40898
rect 0 40840 1858 40896
rect 1914 40840 1919 40896
rect 0 40838 1919 40840
rect 0 40808 800 40838
rect 1853 40835 1919 40838
rect 47301 40898 47367 40901
rect 49200 40898 50000 40928
rect 47301 40896 50000 40898
rect 47301 40840 47306 40896
rect 47362 40840 50000 40896
rect 47301 40838 50000 40840
rect 47301 40835 47367 40838
rect 4208 40832 4528 40833
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 40767 4528 40768
rect 34928 40832 35248 40833
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 49200 40808 50000 40838
rect 34928 40767 35248 40768
rect 20253 40762 20319 40765
rect 20253 40760 20362 40762
rect 20253 40704 20258 40760
rect 20314 40704 20362 40760
rect 20253 40699 20362 40704
rect 20302 40493 20362 40699
rect 20302 40488 20411 40493
rect 20302 40432 20350 40488
rect 20406 40432 20411 40488
rect 20302 40430 20411 40432
rect 20345 40427 20411 40430
rect 19568 40288 19888 40289
rect 0 40218 800 40248
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 40223 19888 40224
rect 1393 40218 1459 40221
rect 0 40216 1459 40218
rect 0 40160 1398 40216
rect 1454 40160 1459 40216
rect 0 40158 1459 40160
rect 0 40128 800 40158
rect 1393 40155 1459 40158
rect 48129 40218 48195 40221
rect 49200 40218 50000 40248
rect 48129 40216 50000 40218
rect 48129 40160 48134 40216
rect 48190 40160 50000 40216
rect 48129 40158 50000 40160
rect 48129 40155 48195 40158
rect 49200 40128 50000 40158
rect 4208 39744 4528 39745
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 39679 4528 39680
rect 34928 39744 35248 39745
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 39679 35248 39680
rect 0 39538 800 39568
rect 2865 39538 2931 39541
rect 0 39536 2931 39538
rect 0 39480 2870 39536
rect 2926 39480 2931 39536
rect 0 39478 2931 39480
rect 0 39448 800 39478
rect 2865 39475 2931 39478
rect 48221 39538 48287 39541
rect 49200 39538 50000 39568
rect 48221 39536 50000 39538
rect 48221 39480 48226 39536
rect 48282 39480 50000 39536
rect 48221 39478 50000 39480
rect 48221 39475 48287 39478
rect 49200 39448 50000 39478
rect 20713 39402 20779 39405
rect 26601 39402 26667 39405
rect 20713 39400 26667 39402
rect 20713 39344 20718 39400
rect 20774 39344 26606 39400
rect 26662 39344 26667 39400
rect 20713 39342 26667 39344
rect 20713 39339 20779 39342
rect 26601 39339 26667 39342
rect 19568 39200 19888 39201
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 39135 19888 39136
rect 0 38768 800 38888
rect 20437 38858 20503 38861
rect 20897 38858 20963 38861
rect 22277 38858 22343 38861
rect 20437 38856 22343 38858
rect 20437 38800 20442 38856
rect 20498 38800 20902 38856
rect 20958 38800 22282 38856
rect 22338 38800 22343 38856
rect 20437 38798 22343 38800
rect 20437 38795 20503 38798
rect 20897 38795 20963 38798
rect 22277 38795 22343 38798
rect 47945 38858 48011 38861
rect 49200 38858 50000 38888
rect 47945 38856 50000 38858
rect 47945 38800 47950 38856
rect 48006 38800 50000 38856
rect 47945 38798 50000 38800
rect 47945 38795 48011 38798
rect 49200 38768 50000 38798
rect 4208 38656 4528 38657
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 38591 4528 38592
rect 34928 38656 35248 38657
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 38591 35248 38592
rect 0 38178 800 38208
rect 4061 38178 4127 38181
rect 0 38176 4127 38178
rect 0 38120 4066 38176
rect 4122 38120 4127 38176
rect 0 38118 4127 38120
rect 0 38088 800 38118
rect 4061 38115 4127 38118
rect 47853 38178 47919 38181
rect 49200 38178 50000 38208
rect 47853 38176 50000 38178
rect 47853 38120 47858 38176
rect 47914 38120 50000 38176
rect 47853 38118 50000 38120
rect 47853 38115 47919 38118
rect 19568 38112 19888 38113
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 49200 38088 50000 38118
rect 19568 38047 19888 38048
rect 4208 37568 4528 37569
rect 0 37498 800 37528
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 1853 37498 1919 37501
rect 0 37496 1919 37498
rect 0 37440 1858 37496
rect 1914 37440 1919 37496
rect 0 37438 1919 37440
rect 0 37408 800 37438
rect 1853 37435 1919 37438
rect 46841 37498 46907 37501
rect 49200 37498 50000 37528
rect 46841 37496 50000 37498
rect 46841 37440 46846 37496
rect 46902 37440 50000 37496
rect 46841 37438 50000 37440
rect 46841 37435 46907 37438
rect 49200 37408 50000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 0 36818 800 36848
rect 1393 36818 1459 36821
rect 0 36816 1459 36818
rect 0 36760 1398 36816
rect 1454 36760 1459 36816
rect 0 36758 1459 36760
rect 0 36728 800 36758
rect 1393 36755 1459 36758
rect 48129 36818 48195 36821
rect 49200 36818 50000 36848
rect 48129 36816 50000 36818
rect 48129 36760 48134 36816
rect 48190 36760 50000 36816
rect 48129 36758 50000 36760
rect 48129 36755 48195 36758
rect 49200 36728 50000 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 2773 36138 2839 36141
rect 0 36136 2839 36138
rect 0 36080 2778 36136
rect 2834 36080 2839 36136
rect 0 36078 2839 36080
rect 0 36048 800 36078
rect 2773 36075 2839 36078
rect 22369 36138 22435 36141
rect 27521 36138 27587 36141
rect 22369 36136 27587 36138
rect 22369 36080 22374 36136
rect 22430 36080 27526 36136
rect 27582 36080 27587 36136
rect 22369 36078 27587 36080
rect 22369 36075 22435 36078
rect 27521 36075 27587 36078
rect 47853 36138 47919 36141
rect 49200 36138 50000 36168
rect 47853 36136 50000 36138
rect 47853 36080 47858 36136
rect 47914 36080 50000 36136
rect 47853 36078 50000 36080
rect 47853 36075 47919 36078
rect 49200 36048 50000 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 20713 35730 20779 35733
rect 21909 35730 21975 35733
rect 20713 35728 21975 35730
rect 20713 35672 20718 35728
rect 20774 35672 21914 35728
rect 21970 35672 21975 35728
rect 20713 35670 21975 35672
rect 20713 35667 20779 35670
rect 21909 35667 21975 35670
rect 26233 35594 26299 35597
rect 27613 35594 27679 35597
rect 26233 35592 27679 35594
rect 26233 35536 26238 35592
rect 26294 35536 27618 35592
rect 27674 35536 27679 35592
rect 26233 35534 27679 35536
rect 26233 35531 26299 35534
rect 27613 35531 27679 35534
rect 0 35368 800 35488
rect 19793 35458 19859 35461
rect 22001 35458 22067 35461
rect 19793 35456 22067 35458
rect 19793 35400 19798 35456
rect 19854 35400 22006 35456
rect 22062 35400 22067 35456
rect 19793 35398 22067 35400
rect 19793 35395 19859 35398
rect 22001 35395 22067 35398
rect 48129 35458 48195 35461
rect 49200 35458 50000 35488
rect 48129 35456 50000 35458
rect 48129 35400 48134 35456
rect 48190 35400 50000 35456
rect 48129 35398 50000 35400
rect 48129 35395 48195 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 49200 35368 50000 35398
rect 34928 35327 35248 35328
rect 19609 35186 19675 35189
rect 24577 35186 24643 35189
rect 19609 35184 24643 35186
rect 19609 35128 19614 35184
rect 19670 35128 24582 35184
rect 24638 35128 24643 35184
rect 19609 35126 24643 35128
rect 19609 35123 19675 35126
rect 24577 35123 24643 35126
rect 19885 35050 19951 35053
rect 21449 35050 21515 35053
rect 21909 35050 21975 35053
rect 19885 35048 21975 35050
rect 19885 34992 19890 35048
rect 19946 34992 21454 35048
rect 21510 34992 21914 35048
rect 21970 34992 21975 35048
rect 19885 34990 21975 34992
rect 19885 34987 19951 34990
rect 21449 34987 21515 34990
rect 21909 34987 21975 34990
rect 19568 34848 19888 34849
rect 0 34778 800 34808
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 1393 34778 1459 34781
rect 0 34776 1459 34778
rect 0 34720 1398 34776
rect 1454 34720 1459 34776
rect 0 34718 1459 34720
rect 0 34688 800 34718
rect 1393 34715 1459 34718
rect 48129 34778 48195 34781
rect 49200 34778 50000 34808
rect 48129 34776 50000 34778
rect 48129 34720 48134 34776
rect 48190 34720 50000 34776
rect 48129 34718 50000 34720
rect 48129 34715 48195 34718
rect 49200 34688 50000 34718
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 0 34098 800 34128
rect 2773 34098 2839 34101
rect 0 34096 2839 34098
rect 0 34040 2778 34096
rect 2834 34040 2839 34096
rect 0 34038 2839 34040
rect 0 34008 800 34038
rect 2773 34035 2839 34038
rect 48037 34098 48103 34101
rect 49200 34098 50000 34128
rect 48037 34096 50000 34098
rect 48037 34040 48042 34096
rect 48098 34040 50000 34096
rect 48037 34038 50000 34040
rect 48037 34035 48103 34038
rect 49200 34008 50000 34038
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 22369 33554 22435 33557
rect 24025 33554 24091 33557
rect 22369 33552 24091 33554
rect 22369 33496 22374 33552
rect 22430 33496 24030 33552
rect 24086 33496 24091 33552
rect 22369 33494 24091 33496
rect 22369 33491 22435 33494
rect 24025 33491 24091 33494
rect 25405 33554 25471 33557
rect 27153 33554 27219 33557
rect 25405 33552 27219 33554
rect 25405 33496 25410 33552
rect 25466 33496 27158 33552
rect 27214 33496 27219 33552
rect 25405 33494 27219 33496
rect 25405 33491 25471 33494
rect 27153 33491 27219 33494
rect 0 33418 800 33448
rect 2773 33418 2839 33421
rect 0 33416 2839 33418
rect 0 33360 2778 33416
rect 2834 33360 2839 33416
rect 0 33358 2839 33360
rect 0 33328 800 33358
rect 2773 33355 2839 33358
rect 47945 33418 48011 33421
rect 49200 33418 50000 33448
rect 47945 33416 50000 33418
rect 47945 33360 47950 33416
rect 48006 33360 50000 33416
rect 47945 33358 50000 33360
rect 47945 33355 48011 33358
rect 49200 33328 50000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 20161 33012 20227 33013
rect 20110 33010 20116 33012
rect 20070 32950 20116 33010
rect 20180 33008 20227 33012
rect 20222 32952 20227 33008
rect 20110 32948 20116 32950
rect 20180 32948 20227 32952
rect 20161 32947 20227 32948
rect 0 32738 800 32768
rect 3141 32738 3207 32741
rect 0 32736 3207 32738
rect 0 32680 3146 32736
rect 3202 32680 3207 32736
rect 0 32678 3207 32680
rect 0 32648 800 32678
rect 3141 32675 3207 32678
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 49200 32648 50000 32768
rect 19568 32607 19888 32608
rect 4208 32128 4528 32129
rect 0 32058 800 32088
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 3233 32058 3299 32061
rect 0 32056 3299 32058
rect 0 32000 3238 32056
rect 3294 32000 3299 32056
rect 0 31998 3299 32000
rect 0 31968 800 31998
rect 3233 31995 3299 31998
rect 47485 32058 47551 32061
rect 49200 32058 50000 32088
rect 47485 32056 50000 32058
rect 47485 32000 47490 32056
rect 47546 32000 50000 32056
rect 47485 31998 50000 32000
rect 47485 31995 47551 31998
rect 49200 31968 50000 31998
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 0 31378 800 31408
rect 1485 31378 1551 31381
rect 0 31376 1551 31378
rect 0 31320 1490 31376
rect 1546 31320 1551 31376
rect 0 31318 1551 31320
rect 0 31288 800 31318
rect 1485 31315 1551 31318
rect 12985 31378 13051 31381
rect 14089 31378 14155 31381
rect 12985 31376 14155 31378
rect 12985 31320 12990 31376
rect 13046 31320 14094 31376
rect 14150 31320 14155 31376
rect 12985 31318 14155 31320
rect 12985 31315 13051 31318
rect 14089 31315 14155 31318
rect 47945 31378 48011 31381
rect 49200 31378 50000 31408
rect 47945 31376 50000 31378
rect 47945 31320 47950 31376
rect 48006 31320 50000 31376
rect 47945 31318 50000 31320
rect 47945 31315 48011 31318
rect 49200 31288 50000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 20253 30834 20319 30837
rect 25773 30834 25839 30837
rect 20253 30832 25839 30834
rect 20253 30776 20258 30832
rect 20314 30776 25778 30832
rect 25834 30776 25839 30832
rect 20253 30774 25839 30776
rect 20253 30771 20319 30774
rect 25773 30771 25839 30774
rect 0 30608 800 30728
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 21081 30290 21147 30293
rect 23422 30290 23428 30292
rect 21081 30288 23428 30290
rect 21081 30232 21086 30288
rect 21142 30232 23428 30288
rect 21081 30230 23428 30232
rect 21081 30227 21147 30230
rect 23422 30228 23428 30230
rect 23492 30228 23498 30292
rect 29269 30290 29335 30293
rect 33225 30290 33291 30293
rect 29269 30288 33291 30290
rect 29269 30232 29274 30288
rect 29330 30232 33230 30288
rect 33286 30232 33291 30288
rect 29269 30230 33291 30232
rect 29269 30227 29335 30230
rect 33225 30227 33291 30230
rect 0 30018 800 30048
rect 2773 30018 2839 30021
rect 0 30016 2839 30018
rect 0 29960 2778 30016
rect 2834 29960 2839 30016
rect 0 29958 2839 29960
rect 0 29928 800 29958
rect 2773 29955 2839 29958
rect 47301 30018 47367 30021
rect 49200 30018 50000 30048
rect 47301 30016 50000 30018
rect 47301 29960 47306 30016
rect 47362 29960 50000 30016
rect 47301 29958 50000 29960
rect 47301 29955 47367 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 49200 29928 50000 29958
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 0 29338 800 29368
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 4061 29338 4127 29341
rect 0 29336 4127 29338
rect 0 29280 4066 29336
rect 4122 29280 4127 29336
rect 0 29278 4127 29280
rect 0 29248 800 29278
rect 4061 29275 4127 29278
rect 46841 29338 46907 29341
rect 49200 29338 50000 29368
rect 46841 29336 50000 29338
rect 46841 29280 46846 29336
rect 46902 29280 50000 29336
rect 46841 29278 50000 29280
rect 46841 29275 46907 29278
rect 49200 29248 50000 29278
rect 19517 29202 19583 29205
rect 20110 29202 20116 29204
rect 19517 29200 20116 29202
rect 19517 29144 19522 29200
rect 19578 29144 20116 29200
rect 19517 29142 20116 29144
rect 19517 29139 19583 29142
rect 20110 29140 20116 29142
rect 20180 29140 20186 29204
rect 16021 29066 16087 29069
rect 18045 29066 18111 29069
rect 16021 29064 18111 29066
rect 16021 29008 16026 29064
rect 16082 29008 18050 29064
rect 18106 29008 18111 29064
rect 16021 29006 18111 29008
rect 16021 29003 16087 29006
rect 18045 29003 18111 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 11145 28794 11211 28797
rect 15653 28794 15719 28797
rect 16757 28794 16823 28797
rect 11145 28792 16823 28794
rect 11145 28736 11150 28792
rect 11206 28736 15658 28792
rect 15714 28736 16762 28792
rect 16818 28736 16823 28792
rect 11145 28734 16823 28736
rect 11145 28731 11211 28734
rect 15653 28731 15719 28734
rect 16757 28731 16823 28734
rect 0 28658 800 28688
rect 2773 28658 2839 28661
rect 0 28656 2839 28658
rect 0 28600 2778 28656
rect 2834 28600 2839 28656
rect 0 28598 2839 28600
rect 0 28568 800 28598
rect 2773 28595 2839 28598
rect 13905 28658 13971 28661
rect 18137 28658 18203 28661
rect 13905 28656 18203 28658
rect 13905 28600 13910 28656
rect 13966 28600 18142 28656
rect 18198 28600 18203 28656
rect 13905 28598 18203 28600
rect 13905 28595 13971 28598
rect 18137 28595 18203 28598
rect 48129 28658 48195 28661
rect 49200 28658 50000 28688
rect 48129 28656 50000 28658
rect 48129 28600 48134 28656
rect 48190 28600 50000 28656
rect 48129 28598 50000 28600
rect 48129 28595 48195 28598
rect 49200 28568 50000 28598
rect 12065 28522 12131 28525
rect 17677 28522 17743 28525
rect 12065 28520 17743 28522
rect 12065 28464 12070 28520
rect 12126 28464 17682 28520
rect 17738 28464 17743 28520
rect 12065 28462 17743 28464
rect 12065 28459 12131 28462
rect 17677 28459 17743 28462
rect 20805 28386 20871 28389
rect 27889 28386 27955 28389
rect 20805 28384 27955 28386
rect 20805 28328 20810 28384
rect 20866 28328 27894 28384
rect 27950 28328 27955 28384
rect 20805 28326 27955 28328
rect 20805 28323 20871 28326
rect 27889 28323 27955 28326
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 27429 28114 27495 28117
rect 28073 28114 28139 28117
rect 29269 28114 29335 28117
rect 27429 28112 29335 28114
rect 27429 28056 27434 28112
rect 27490 28056 28078 28112
rect 28134 28056 29274 28112
rect 29330 28056 29335 28112
rect 27429 28054 29335 28056
rect 27429 28051 27495 28054
rect 28073 28051 28139 28054
rect 29269 28051 29335 28054
rect 0 27888 800 28008
rect 47853 27978 47919 27981
rect 49200 27978 50000 28008
rect 47853 27976 50000 27978
rect 47853 27920 47858 27976
rect 47914 27920 50000 27976
rect 47853 27918 50000 27920
rect 47853 27915 47919 27918
rect 49200 27888 50000 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 19701 27434 19767 27437
rect 20069 27434 20135 27437
rect 19701 27432 20135 27434
rect 19701 27376 19706 27432
rect 19762 27376 20074 27432
rect 20130 27376 20135 27432
rect 19701 27374 20135 27376
rect 19701 27371 19767 27374
rect 20069 27371 20135 27374
rect 0 27298 800 27328
rect 2773 27298 2839 27301
rect 0 27296 2839 27298
rect 0 27240 2778 27296
rect 2834 27240 2839 27296
rect 0 27238 2839 27240
rect 0 27208 800 27238
rect 2773 27235 2839 27238
rect 23749 27298 23815 27301
rect 27981 27298 28047 27301
rect 28625 27298 28691 27301
rect 23749 27296 28691 27298
rect 23749 27240 23754 27296
rect 23810 27240 27986 27296
rect 28042 27240 28630 27296
rect 28686 27240 28691 27296
rect 23749 27238 28691 27240
rect 23749 27235 23815 27238
rect 27981 27235 28047 27238
rect 28625 27235 28691 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 49200 27208 50000 27328
rect 19568 27167 19888 27168
rect 23381 27026 23447 27029
rect 27429 27026 27495 27029
rect 23381 27024 27495 27026
rect 23381 26968 23386 27024
rect 23442 26968 27434 27024
rect 27490 26968 27495 27024
rect 23381 26966 27495 26968
rect 23381 26963 23447 26966
rect 27429 26963 27495 26966
rect 29545 26754 29611 26757
rect 32397 26754 32463 26757
rect 29545 26752 32463 26754
rect 29545 26696 29550 26752
rect 29606 26696 32402 26752
rect 32458 26696 32463 26752
rect 29545 26694 32463 26696
rect 29545 26691 29611 26694
rect 32397 26691 32463 26694
rect 4208 26688 4528 26689
rect 0 26618 800 26648
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 2773 26618 2839 26621
rect 0 26616 2839 26618
rect 0 26560 2778 26616
rect 2834 26560 2839 26616
rect 0 26558 2839 26560
rect 0 26528 800 26558
rect 2773 26555 2839 26558
rect 45553 26618 45619 26621
rect 49200 26618 50000 26648
rect 45553 26616 50000 26618
rect 45553 26560 45558 26616
rect 45614 26560 50000 26616
rect 45553 26558 50000 26560
rect 45553 26555 45619 26558
rect 49200 26528 50000 26558
rect 15469 26346 15535 26349
rect 17677 26346 17743 26349
rect 15469 26344 17743 26346
rect 15469 26288 15474 26344
rect 15530 26288 17682 26344
rect 17738 26288 17743 26344
rect 15469 26286 17743 26288
rect 15469 26283 15535 26286
rect 17677 26283 17743 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 0 25938 800 25968
rect 1577 25938 1643 25941
rect 0 25936 1643 25938
rect 0 25880 1582 25936
rect 1638 25880 1643 25936
rect 0 25878 1643 25880
rect 0 25848 800 25878
rect 1577 25875 1643 25878
rect 12709 25938 12775 25941
rect 17401 25938 17467 25941
rect 12709 25936 17467 25938
rect 12709 25880 12714 25936
rect 12770 25880 17406 25936
rect 17462 25880 17467 25936
rect 12709 25878 17467 25880
rect 12709 25875 12775 25878
rect 17401 25875 17467 25878
rect 47945 25938 48011 25941
rect 49200 25938 50000 25968
rect 47945 25936 50000 25938
rect 47945 25880 47950 25936
rect 48006 25880 50000 25936
rect 47945 25878 50000 25880
rect 47945 25875 48011 25878
rect 49200 25848 50000 25878
rect 14273 25802 14339 25805
rect 17125 25802 17191 25805
rect 14273 25800 17191 25802
rect 14273 25744 14278 25800
rect 14334 25744 17130 25800
rect 17186 25744 17191 25800
rect 14273 25742 17191 25744
rect 14273 25739 14339 25742
rect 17125 25739 17191 25742
rect 16205 25666 16271 25669
rect 18229 25666 18295 25669
rect 16205 25664 18295 25666
rect 16205 25608 16210 25664
rect 16266 25608 18234 25664
rect 18290 25608 18295 25664
rect 16205 25606 18295 25608
rect 16205 25603 16271 25606
rect 18229 25603 18295 25606
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 0 25168 800 25288
rect 47853 25258 47919 25261
rect 49200 25258 50000 25288
rect 47853 25256 50000 25258
rect 47853 25200 47858 25256
rect 47914 25200 50000 25256
rect 47853 25198 50000 25200
rect 47853 25195 47919 25198
rect 49200 25168 50000 25198
rect 23105 25122 23171 25125
rect 24342 25122 24348 25124
rect 23105 25120 24348 25122
rect 23105 25064 23110 25120
rect 23166 25064 24348 25120
rect 23105 25062 24348 25064
rect 23105 25059 23171 25062
rect 24342 25060 24348 25062
rect 24412 25122 24418 25124
rect 24485 25122 24551 25125
rect 24412 25120 24551 25122
rect 24412 25064 24490 25120
rect 24546 25064 24551 25120
rect 24412 25062 24551 25064
rect 24412 25060 24418 25062
rect 24485 25059 24551 25062
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 20069 24986 20135 24989
rect 24669 24986 24735 24989
rect 27153 24986 27219 24989
rect 20069 24984 27219 24986
rect 20069 24928 20074 24984
rect 20130 24928 24674 24984
rect 24730 24928 27158 24984
rect 27214 24928 27219 24984
rect 20069 24926 27219 24928
rect 20069 24923 20135 24926
rect 24669 24923 24735 24926
rect 27153 24923 27219 24926
rect 20345 24850 20411 24853
rect 38101 24850 38167 24853
rect 20345 24848 38167 24850
rect 20345 24792 20350 24848
rect 20406 24792 38106 24848
rect 38162 24792 38167 24848
rect 20345 24790 38167 24792
rect 20345 24787 20411 24790
rect 38101 24787 38167 24790
rect 19977 24714 20043 24717
rect 21357 24714 21423 24717
rect 19977 24712 21423 24714
rect 19977 24656 19982 24712
rect 20038 24656 21362 24712
rect 21418 24656 21423 24712
rect 19977 24654 21423 24656
rect 19977 24651 20043 24654
rect 21357 24651 21423 24654
rect 0 24488 800 24608
rect 20345 24578 20411 24581
rect 21633 24578 21699 24581
rect 20345 24576 21699 24578
rect 20345 24520 20350 24576
rect 20406 24520 21638 24576
rect 21694 24520 21699 24576
rect 20345 24518 21699 24520
rect 20345 24515 20411 24518
rect 21633 24515 21699 24518
rect 22921 24578 22987 24581
rect 24209 24578 24275 24581
rect 25865 24578 25931 24581
rect 22921 24576 25931 24578
rect 22921 24520 22926 24576
rect 22982 24520 24214 24576
rect 24270 24520 25870 24576
rect 25926 24520 25931 24576
rect 22921 24518 25931 24520
rect 22921 24515 22987 24518
rect 24209 24515 24275 24518
rect 25865 24515 25931 24518
rect 48129 24578 48195 24581
rect 49200 24578 50000 24608
rect 48129 24576 50000 24578
rect 48129 24520 48134 24576
rect 48190 24520 50000 24576
rect 48129 24518 50000 24520
rect 48129 24515 48195 24518
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 49200 24488 50000 24518
rect 34928 24447 35248 24448
rect 20069 24442 20135 24445
rect 21173 24442 21239 24445
rect 20069 24440 21239 24442
rect 20069 24384 20074 24440
rect 20130 24384 21178 24440
rect 21234 24384 21239 24440
rect 20069 24382 21239 24384
rect 20069 24379 20135 24382
rect 21173 24379 21239 24382
rect 19885 24306 19951 24309
rect 26601 24306 26667 24309
rect 19885 24304 26667 24306
rect 19885 24248 19890 24304
rect 19946 24248 26606 24304
rect 26662 24248 26667 24304
rect 19885 24246 26667 24248
rect 19885 24243 19951 24246
rect 26601 24243 26667 24246
rect 23841 24170 23907 24173
rect 24669 24170 24735 24173
rect 23841 24168 24735 24170
rect 23841 24112 23846 24168
rect 23902 24112 24674 24168
rect 24730 24112 24735 24168
rect 23841 24110 24735 24112
rect 23841 24107 23907 24110
rect 24669 24107 24735 24110
rect 24577 24034 24643 24037
rect 28901 24034 28967 24037
rect 24577 24032 28967 24034
rect 24577 23976 24582 24032
rect 24638 23976 28906 24032
rect 28962 23976 28967 24032
rect 24577 23974 28967 23976
rect 24577 23971 24643 23974
rect 28901 23971 28967 23974
rect 19568 23968 19888 23969
rect 0 23898 800 23928
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 1393 23898 1459 23901
rect 0 23896 1459 23898
rect 0 23840 1398 23896
rect 1454 23840 1459 23896
rect 0 23838 1459 23840
rect 0 23808 800 23838
rect 1393 23835 1459 23838
rect 47945 23898 48011 23901
rect 49200 23898 50000 23928
rect 47945 23896 50000 23898
rect 47945 23840 47950 23896
rect 48006 23840 50000 23896
rect 47945 23838 50000 23840
rect 47945 23835 48011 23838
rect 49200 23808 50000 23838
rect 18045 23762 18111 23765
rect 47577 23762 47643 23765
rect 18045 23760 47643 23762
rect 18045 23704 18050 23760
rect 18106 23704 47582 23760
rect 47638 23704 47643 23760
rect 18045 23702 47643 23704
rect 18045 23699 18111 23702
rect 47577 23699 47643 23702
rect 11973 23626 12039 23629
rect 18413 23626 18479 23629
rect 11973 23624 18479 23626
rect 11973 23568 11978 23624
rect 12034 23568 18418 23624
rect 18474 23568 18479 23624
rect 11973 23566 18479 23568
rect 11973 23563 12039 23566
rect 18413 23563 18479 23566
rect 20345 23626 20411 23629
rect 26233 23626 26299 23629
rect 20345 23624 26299 23626
rect 20345 23568 20350 23624
rect 20406 23568 26238 23624
rect 26294 23568 26299 23624
rect 20345 23566 26299 23568
rect 20345 23563 20411 23566
rect 26233 23563 26299 23566
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 2773 23218 2839 23221
rect 0 23216 2839 23218
rect 0 23160 2778 23216
rect 2834 23160 2839 23216
rect 0 23158 2839 23160
rect 0 23128 800 23158
rect 2773 23155 2839 23158
rect 49200 23128 50000 23248
rect 10317 23082 10383 23085
rect 14457 23082 14523 23085
rect 10317 23080 14523 23082
rect 10317 23024 10322 23080
rect 10378 23024 14462 23080
rect 14518 23024 14523 23080
rect 10317 23022 14523 23024
rect 10317 23019 10383 23022
rect 14457 23019 14523 23022
rect 23422 22884 23428 22948
rect 23492 22946 23498 22948
rect 24393 22946 24459 22949
rect 23492 22944 24459 22946
rect 23492 22888 24398 22944
rect 24454 22888 24459 22944
rect 23492 22886 24459 22888
rect 23492 22884 23498 22886
rect 24393 22883 24459 22886
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 0 22538 800 22568
rect 1853 22538 1919 22541
rect 0 22536 1919 22538
rect 0 22480 1858 22536
rect 1914 22480 1919 22536
rect 0 22478 1919 22480
rect 0 22448 800 22478
rect 1853 22475 1919 22478
rect 17677 22538 17743 22541
rect 23565 22538 23631 22541
rect 17677 22536 23631 22538
rect 17677 22480 17682 22536
rect 17738 22480 23570 22536
rect 23626 22480 23631 22536
rect 17677 22478 23631 22480
rect 17677 22475 17743 22478
rect 23565 22475 23631 22478
rect 48129 22538 48195 22541
rect 49200 22538 50000 22568
rect 48129 22536 50000 22538
rect 48129 22480 48134 22536
rect 48190 22480 50000 22536
rect 48129 22478 50000 22480
rect 48129 22475 48195 22478
rect 49200 22448 50000 22478
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 20253 21994 20319 21997
rect 22093 21994 22159 21997
rect 20253 21992 22159 21994
rect 20253 21936 20258 21992
rect 20314 21936 22098 21992
rect 22154 21936 22159 21992
rect 20253 21934 22159 21936
rect 20253 21931 20319 21934
rect 22093 21931 22159 21934
rect 0 21858 800 21888
rect 3969 21858 4035 21861
rect 0 21856 4035 21858
rect 0 21800 3974 21856
rect 4030 21800 4035 21856
rect 0 21798 4035 21800
rect 0 21768 800 21798
rect 3969 21795 4035 21798
rect 24577 21858 24643 21861
rect 27797 21858 27863 21861
rect 24577 21856 27863 21858
rect 24577 21800 24582 21856
rect 24638 21800 27802 21856
rect 27858 21800 27863 21856
rect 24577 21798 27863 21800
rect 24577 21795 24643 21798
rect 27797 21795 27863 21798
rect 47945 21858 48011 21861
rect 49200 21858 50000 21888
rect 47945 21856 50000 21858
rect 47945 21800 47950 21856
rect 48006 21800 50000 21856
rect 47945 21798 50000 21800
rect 47945 21795 48011 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 49200 21768 50000 21798
rect 19568 21727 19888 21728
rect 20989 21722 21055 21725
rect 24577 21722 24643 21725
rect 20989 21720 24643 21722
rect 20989 21664 20994 21720
rect 21050 21664 24582 21720
rect 24638 21664 24643 21720
rect 20989 21662 24643 21664
rect 20989 21659 21055 21662
rect 24577 21659 24643 21662
rect 20713 21586 20779 21589
rect 21173 21586 21239 21589
rect 20713 21584 21239 21586
rect 20713 21528 20718 21584
rect 20774 21528 21178 21584
rect 21234 21528 21239 21584
rect 20713 21526 21239 21528
rect 20713 21523 20779 21526
rect 21173 21523 21239 21526
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 4061 21178 4127 21181
rect 0 21176 4127 21178
rect 0 21120 4066 21176
rect 4122 21120 4127 21176
rect 0 21118 4127 21120
rect 0 21088 800 21118
rect 4061 21115 4127 21118
rect 49200 21088 50000 21208
rect 24393 20770 24459 20773
rect 24526 20770 24532 20772
rect 24393 20768 24532 20770
rect 24393 20712 24398 20768
rect 24454 20712 24532 20768
rect 24393 20710 24532 20712
rect 24393 20707 24459 20710
rect 24526 20708 24532 20710
rect 24596 20708 24602 20772
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 0 20408 800 20528
rect 10961 20498 11027 20501
rect 12433 20498 12499 20501
rect 10961 20496 12499 20498
rect 10961 20440 10966 20496
rect 11022 20440 12438 20496
rect 12494 20440 12499 20496
rect 10961 20438 12499 20440
rect 10961 20435 11027 20438
rect 12433 20435 12499 20438
rect 23289 20498 23355 20501
rect 24342 20498 24348 20500
rect 23289 20496 24348 20498
rect 23289 20440 23294 20496
rect 23350 20440 24348 20496
rect 23289 20438 24348 20440
rect 23289 20435 23355 20438
rect 24342 20436 24348 20438
rect 24412 20498 24418 20500
rect 26233 20498 26299 20501
rect 24412 20496 26299 20498
rect 24412 20440 26238 20496
rect 26294 20440 26299 20496
rect 24412 20438 26299 20440
rect 24412 20436 24418 20438
rect 26233 20435 26299 20438
rect 49200 20408 50000 20528
rect 15929 20362 15995 20365
rect 18597 20362 18663 20365
rect 15929 20360 18663 20362
rect 15929 20304 15934 20360
rect 15990 20304 18602 20360
rect 18658 20304 18663 20360
rect 15929 20302 18663 20304
rect 15929 20299 15995 20302
rect 18597 20299 18663 20302
rect 23197 20362 23263 20365
rect 23974 20362 23980 20364
rect 23197 20360 23980 20362
rect 23197 20304 23202 20360
rect 23258 20304 23980 20360
rect 23197 20302 23980 20304
rect 23197 20299 23263 20302
rect 23974 20300 23980 20302
rect 24044 20300 24050 20364
rect 12249 20226 12315 20229
rect 17493 20226 17559 20229
rect 12249 20224 17559 20226
rect 12249 20168 12254 20224
rect 12310 20168 17498 20224
rect 17554 20168 17559 20224
rect 12249 20166 17559 20168
rect 12249 20163 12315 20166
rect 17493 20163 17559 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 11973 19954 12039 19957
rect 14273 19954 14339 19957
rect 11973 19952 14339 19954
rect 11973 19896 11978 19952
rect 12034 19896 14278 19952
rect 14334 19896 14339 19952
rect 11973 19894 14339 19896
rect 11973 19891 12039 19894
rect 14273 19891 14339 19894
rect 0 19818 800 19848
rect 4061 19818 4127 19821
rect 0 19816 4127 19818
rect 0 19760 4066 19816
rect 4122 19760 4127 19816
rect 0 19758 4127 19760
rect 0 19728 800 19758
rect 4061 19755 4127 19758
rect 12617 19818 12683 19821
rect 17677 19818 17743 19821
rect 18689 19818 18755 19821
rect 12617 19816 18755 19818
rect 12617 19760 12622 19816
rect 12678 19760 17682 19816
rect 17738 19760 18694 19816
rect 18750 19760 18755 19816
rect 12617 19758 18755 19760
rect 12617 19755 12683 19758
rect 17677 19755 17743 19758
rect 18689 19755 18755 19758
rect 48129 19818 48195 19821
rect 49200 19818 50000 19848
rect 48129 19816 50000 19818
rect 48129 19760 48134 19816
rect 48190 19760 50000 19816
rect 48129 19758 50000 19760
rect 48129 19755 48195 19758
rect 49200 19728 50000 19758
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 11973 19546 12039 19549
rect 13261 19546 13327 19549
rect 11973 19544 13327 19546
rect 11973 19488 11978 19544
rect 12034 19488 13266 19544
rect 13322 19488 13327 19544
rect 11973 19486 13327 19488
rect 11973 19483 12039 19486
rect 13261 19483 13327 19486
rect 18229 19546 18295 19549
rect 19057 19546 19123 19549
rect 18229 19544 19123 19546
rect 18229 19488 18234 19544
rect 18290 19488 19062 19544
rect 19118 19488 19123 19544
rect 18229 19486 19123 19488
rect 18229 19483 18295 19486
rect 19057 19483 19123 19486
rect 25681 19410 25747 19413
rect 25681 19408 25882 19410
rect 25681 19352 25686 19408
rect 25742 19352 25882 19408
rect 25681 19350 25882 19352
rect 25681 19347 25747 19350
rect 25822 19274 25882 19350
rect 26325 19274 26391 19277
rect 25822 19272 26391 19274
rect 25822 19216 26330 19272
rect 26386 19216 26391 19272
rect 25822 19214 26391 19216
rect 26325 19211 26391 19214
rect 0 19138 800 19168
rect 2773 19138 2839 19141
rect 0 19136 2839 19138
rect 0 19080 2778 19136
rect 2834 19080 2839 19136
rect 0 19078 2839 19080
rect 0 19048 800 19078
rect 2773 19075 2839 19078
rect 47301 19138 47367 19141
rect 49200 19138 50000 19168
rect 47301 19136 50000 19138
rect 47301 19080 47306 19136
rect 47362 19080 50000 19136
rect 47301 19078 50000 19080
rect 47301 19075 47367 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 49200 19048 50000 19078
rect 34928 19007 35248 19008
rect 19568 18528 19888 18529
rect 0 18458 800 18488
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 3141 18458 3207 18461
rect 0 18456 3207 18458
rect 0 18400 3146 18456
rect 3202 18400 3207 18456
rect 0 18398 3207 18400
rect 0 18368 800 18398
rect 3141 18395 3207 18398
rect 22093 18458 22159 18461
rect 28165 18458 28231 18461
rect 22093 18456 28231 18458
rect 22093 18400 22098 18456
rect 22154 18400 28170 18456
rect 28226 18400 28231 18456
rect 22093 18398 28231 18400
rect 22093 18395 22159 18398
rect 28165 18395 28231 18398
rect 49200 18368 50000 18488
rect 10961 18322 11027 18325
rect 12249 18322 12315 18325
rect 10961 18320 12315 18322
rect 10961 18264 10966 18320
rect 11022 18264 12254 18320
rect 12310 18264 12315 18320
rect 10961 18262 12315 18264
rect 10961 18259 11027 18262
rect 12249 18259 12315 18262
rect 20621 18322 20687 18325
rect 25313 18322 25379 18325
rect 26049 18322 26115 18325
rect 20621 18320 25379 18322
rect 20621 18264 20626 18320
rect 20682 18264 25318 18320
rect 25374 18264 25379 18320
rect 20621 18262 25379 18264
rect 20621 18259 20687 18262
rect 25313 18259 25379 18262
rect 25822 18320 26115 18322
rect 25822 18264 26054 18320
rect 26110 18264 26115 18320
rect 25822 18262 26115 18264
rect 25681 18186 25747 18189
rect 25822 18186 25882 18262
rect 26049 18259 26115 18262
rect 25681 18184 25882 18186
rect 25681 18128 25686 18184
rect 25742 18128 25882 18184
rect 25681 18126 25882 18128
rect 25681 18123 25747 18126
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 21817 17914 21883 17917
rect 28441 17914 28507 17917
rect 21817 17912 28507 17914
rect 21817 17856 21822 17912
rect 21878 17856 28446 17912
rect 28502 17856 28507 17912
rect 21817 17854 28507 17856
rect 21817 17851 21883 17854
rect 28441 17851 28507 17854
rect 0 17778 800 17808
rect 2773 17778 2839 17781
rect 28165 17780 28231 17781
rect 28165 17778 28212 17780
rect 0 17776 2839 17778
rect 0 17720 2778 17776
rect 2834 17720 2839 17776
rect 0 17718 2839 17720
rect 28120 17776 28212 17778
rect 28120 17720 28170 17776
rect 28120 17718 28212 17720
rect 0 17688 800 17718
rect 2773 17715 2839 17718
rect 28165 17716 28212 17718
rect 28276 17716 28282 17780
rect 45645 17778 45711 17781
rect 49200 17778 50000 17808
rect 45645 17776 50000 17778
rect 45645 17720 45650 17776
rect 45706 17720 50000 17776
rect 45645 17718 50000 17720
rect 28165 17715 28231 17716
rect 45645 17715 45711 17718
rect 49200 17688 50000 17718
rect 23381 17642 23447 17645
rect 23381 17640 23674 17642
rect 23381 17584 23386 17640
rect 23442 17584 23674 17640
rect 23381 17582 23674 17584
rect 23381 17579 23447 17582
rect 20161 17506 20227 17509
rect 22645 17506 22711 17509
rect 23381 17506 23447 17509
rect 20161 17504 20362 17506
rect 20161 17448 20166 17504
rect 20222 17448 20362 17504
rect 20161 17446 20362 17448
rect 20161 17443 20227 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 20302 17373 20362 17446
rect 22645 17504 23447 17506
rect 22645 17448 22650 17504
rect 22706 17448 23386 17504
rect 23442 17448 23447 17504
rect 22645 17446 23447 17448
rect 22645 17443 22711 17446
rect 23381 17443 23447 17446
rect 20302 17368 20411 17373
rect 20302 17312 20350 17368
rect 20406 17312 20411 17368
rect 20302 17310 20411 17312
rect 20345 17307 20411 17310
rect 22921 17370 22987 17373
rect 23614 17370 23674 17582
rect 22921 17368 23674 17370
rect 22921 17312 22926 17368
rect 22982 17312 23674 17368
rect 22921 17310 23674 17312
rect 22921 17307 22987 17310
rect 0 17098 800 17128
rect 1853 17098 1919 17101
rect 0 17096 1919 17098
rect 0 17040 1858 17096
rect 1914 17040 1919 17096
rect 0 17038 1919 17040
rect 0 17008 800 17038
rect 1853 17035 1919 17038
rect 22461 17098 22527 17101
rect 23657 17098 23723 17101
rect 22461 17096 23723 17098
rect 22461 17040 22466 17096
rect 22522 17040 23662 17096
rect 23718 17040 23723 17096
rect 22461 17038 23723 17040
rect 22461 17035 22527 17038
rect 23657 17035 23723 17038
rect 48129 17098 48195 17101
rect 49200 17098 50000 17128
rect 48129 17096 50000 17098
rect 48129 17040 48134 17096
rect 48190 17040 50000 17096
rect 48129 17038 50000 17040
rect 48129 17035 48195 17038
rect 49200 17008 50000 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 23381 16826 23447 16829
rect 44817 16826 44883 16829
rect 45645 16826 45711 16829
rect 23381 16824 23674 16826
rect 23381 16768 23386 16824
rect 23442 16768 23674 16824
rect 23381 16766 23674 16768
rect 23381 16763 23447 16766
rect 22369 16690 22435 16693
rect 23614 16690 23674 16766
rect 44817 16824 45711 16826
rect 44817 16768 44822 16824
rect 44878 16768 45650 16824
rect 45706 16768 45711 16824
rect 44817 16766 45711 16768
rect 44817 16763 44883 16766
rect 45645 16763 45711 16766
rect 23841 16690 23907 16693
rect 22369 16688 23490 16690
rect 22369 16632 22374 16688
rect 22430 16632 23490 16688
rect 22369 16630 23490 16632
rect 23614 16688 23907 16690
rect 23614 16632 23846 16688
rect 23902 16632 23907 16688
rect 23614 16630 23907 16632
rect 22369 16627 22435 16630
rect 23430 16557 23490 16630
rect 23841 16627 23907 16630
rect 23430 16552 23539 16557
rect 23430 16496 23478 16552
rect 23534 16496 23539 16552
rect 23430 16494 23539 16496
rect 23473 16491 23539 16494
rect 0 16418 800 16448
rect 2773 16418 2839 16421
rect 0 16416 2839 16418
rect 0 16360 2778 16416
rect 2834 16360 2839 16416
rect 0 16358 2839 16360
rect 0 16328 800 16358
rect 2773 16355 2839 16358
rect 28206 16356 28212 16420
rect 28276 16418 28282 16420
rect 28349 16418 28415 16421
rect 28276 16416 28415 16418
rect 28276 16360 28354 16416
rect 28410 16360 28415 16416
rect 28276 16358 28415 16360
rect 28276 16356 28282 16358
rect 28349 16355 28415 16358
rect 48129 16418 48195 16421
rect 49200 16418 50000 16448
rect 48129 16416 50000 16418
rect 48129 16360 48134 16416
rect 48190 16360 50000 16416
rect 48129 16358 50000 16360
rect 48129 16355 48195 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 49200 16328 50000 16358
rect 19568 16287 19888 16288
rect 22921 16146 22987 16149
rect 23657 16146 23723 16149
rect 26141 16146 26207 16149
rect 22921 16144 26207 16146
rect 22921 16088 22926 16144
rect 22982 16088 23662 16144
rect 23718 16088 26146 16144
rect 26202 16088 26207 16144
rect 22921 16086 26207 16088
rect 22921 16083 22987 16086
rect 23657 16083 23723 16086
rect 26141 16083 26207 16086
rect 30005 16010 30071 16013
rect 30281 16010 30347 16013
rect 31017 16010 31083 16013
rect 30005 16008 31083 16010
rect 30005 15952 30010 16008
rect 30066 15952 30286 16008
rect 30342 15952 31022 16008
rect 31078 15952 31083 16008
rect 30005 15950 31083 15952
rect 30005 15947 30071 15950
rect 30281 15947 30347 15950
rect 31017 15947 31083 15950
rect 29545 15874 29611 15877
rect 32305 15874 32371 15877
rect 29545 15872 32371 15874
rect 29545 15816 29550 15872
rect 29606 15816 32310 15872
rect 32366 15816 32371 15872
rect 29545 15814 32371 15816
rect 29545 15811 29611 15814
rect 32305 15811 32371 15814
rect 4208 15808 4528 15809
rect 0 15648 800 15768
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 27613 15738 27679 15741
rect 27797 15738 27863 15741
rect 30741 15738 30807 15741
rect 27613 15736 30807 15738
rect 27613 15680 27618 15736
rect 27674 15680 27802 15736
rect 27858 15680 30746 15736
rect 30802 15680 30807 15736
rect 27613 15678 30807 15680
rect 27613 15675 27679 15678
rect 27797 15675 27863 15678
rect 30741 15675 30807 15678
rect 49200 15648 50000 15768
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 0 14968 800 15088
rect 46841 15058 46907 15061
rect 49200 15058 50000 15088
rect 46841 15056 50000 15058
rect 46841 15000 46846 15056
rect 46902 15000 50000 15056
rect 46841 14998 50000 15000
rect 46841 14995 46907 14998
rect 49200 14968 50000 14998
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14288 800 14408
rect 48129 14378 48195 14381
rect 49200 14378 50000 14408
rect 48129 14376 50000 14378
rect 48129 14320 48134 14376
rect 48190 14320 50000 14376
rect 48129 14318 50000 14320
rect 48129 14315 48195 14318
rect 49200 14288 50000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 0 13698 800 13728
rect 2773 13698 2839 13701
rect 0 13696 2839 13698
rect 0 13640 2778 13696
rect 2834 13640 2839 13696
rect 0 13638 2839 13640
rect 0 13608 800 13638
rect 2773 13635 2839 13638
rect 47853 13698 47919 13701
rect 49200 13698 50000 13728
rect 47853 13696 50000 13698
rect 47853 13640 47858 13696
rect 47914 13640 50000 13696
rect 47853 13638 50000 13640
rect 47853 13635 47919 13638
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 49200 13608 50000 13638
rect 34928 13567 35248 13568
rect 19568 13088 19888 13089
rect 0 13018 800 13048
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 4061 13018 4127 13021
rect 0 13016 4127 13018
rect 0 12960 4066 13016
rect 4122 12960 4127 13016
rect 0 12958 4127 12960
rect 0 12928 800 12958
rect 4061 12955 4127 12958
rect 46841 13018 46907 13021
rect 49200 13018 50000 13048
rect 46841 13016 50000 13018
rect 46841 12960 46846 13016
rect 46902 12960 50000 13016
rect 46841 12958 50000 12960
rect 46841 12955 46907 12958
rect 49200 12928 50000 12958
rect 26233 12746 26299 12749
rect 27245 12746 27311 12749
rect 26233 12744 27311 12746
rect 26233 12688 26238 12744
rect 26294 12688 27250 12744
rect 27306 12688 27311 12744
rect 26233 12686 27311 12688
rect 26233 12683 26299 12686
rect 27245 12683 27311 12686
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 45553 12338 45619 12341
rect 49200 12338 50000 12368
rect 45553 12336 50000 12338
rect 45553 12280 45558 12336
rect 45614 12280 50000 12336
rect 45553 12278 50000 12280
rect 45553 12275 45619 12278
rect 49200 12248 50000 12278
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 0 11568 800 11688
rect 49200 11568 50000 11688
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 28993 11114 29059 11117
rect 28950 11112 29059 11114
rect 28950 11056 28998 11112
rect 29054 11056 29059 11112
rect 28950 11051 29059 11056
rect 0 10978 800 11008
rect 1393 10978 1459 10981
rect 0 10976 1459 10978
rect 0 10920 1398 10976
rect 1454 10920 1459 10976
rect 0 10918 1459 10920
rect 0 10888 800 10918
rect 1393 10915 1459 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 28950 10437 29010 11051
rect 48129 10978 48195 10981
rect 49200 10978 50000 11008
rect 48129 10976 50000 10978
rect 48129 10920 48134 10976
rect 48190 10920 50000 10976
rect 48129 10918 50000 10920
rect 48129 10915 48195 10918
rect 49200 10888 50000 10918
rect 28950 10432 29059 10437
rect 28950 10376 28998 10432
rect 29054 10376 29059 10432
rect 28950 10374 29059 10376
rect 28993 10371 29059 10374
rect 29361 10434 29427 10437
rect 30925 10434 30991 10437
rect 29361 10432 30991 10434
rect 29361 10376 29366 10432
rect 29422 10376 30930 10432
rect 30986 10376 30991 10432
rect 29361 10374 30991 10376
rect 29361 10371 29427 10374
rect 30925 10371 30991 10374
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 3049 10298 3115 10301
rect 0 10296 3115 10298
rect 0 10240 3054 10296
rect 3110 10240 3115 10296
rect 0 10238 3115 10240
rect 0 10208 800 10238
rect 3049 10235 3115 10238
rect 47761 10298 47827 10301
rect 49200 10298 50000 10328
rect 47761 10296 50000 10298
rect 47761 10240 47766 10296
rect 47822 10240 50000 10296
rect 47761 10238 50000 10240
rect 47761 10235 47827 10238
rect 49200 10208 50000 10238
rect 26785 10026 26851 10029
rect 28901 10026 28967 10029
rect 26785 10024 28967 10026
rect 26785 9968 26790 10024
rect 26846 9968 28906 10024
rect 28962 9968 28967 10024
rect 26785 9966 28967 9968
rect 26785 9963 26851 9966
rect 28901 9963 28967 9966
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 0 9618 800 9648
rect 3233 9618 3299 9621
rect 0 9616 3299 9618
rect 0 9560 3238 9616
rect 3294 9560 3299 9616
rect 0 9558 3299 9560
rect 0 9528 800 9558
rect 3233 9555 3299 9558
rect 46381 9618 46447 9621
rect 49200 9618 50000 9648
rect 46381 9616 50000 9618
rect 46381 9560 46386 9616
rect 46442 9560 50000 9616
rect 46381 9558 50000 9560
rect 46381 9555 46447 9558
rect 49200 9528 50000 9558
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 0 8938 800 8968
rect 2957 8938 3023 8941
rect 0 8936 3023 8938
rect 0 8880 2962 8936
rect 3018 8880 3023 8936
rect 0 8878 3023 8880
rect 0 8848 800 8878
rect 2957 8875 3023 8878
rect 47945 8938 48011 8941
rect 49200 8938 50000 8968
rect 47945 8936 50000 8938
rect 47945 8880 47950 8936
rect 48006 8880 50000 8936
rect 47945 8878 50000 8880
rect 47945 8875 48011 8878
rect 49200 8848 50000 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 0 8258 800 8288
rect 1853 8258 1919 8261
rect 0 8256 1919 8258
rect 0 8200 1858 8256
rect 1914 8200 1919 8256
rect 0 8198 1919 8200
rect 0 8168 800 8198
rect 1853 8195 1919 8198
rect 47761 8258 47827 8261
rect 49200 8258 50000 8288
rect 47761 8256 50000 8258
rect 47761 8200 47766 8256
rect 47822 8200 50000 8256
rect 47761 8198 50000 8200
rect 47761 8195 47827 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 49200 8168 50000 8198
rect 34928 8127 35248 8128
rect 19568 7648 19888 7649
rect 0 7578 800 7608
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 1853 7578 1919 7581
rect 0 7576 1919 7578
rect 0 7520 1858 7576
rect 1914 7520 1919 7576
rect 0 7518 1919 7520
rect 0 7488 800 7518
rect 1853 7515 1919 7518
rect 48129 7578 48195 7581
rect 49200 7578 50000 7608
rect 48129 7576 50000 7578
rect 48129 7520 48134 7576
rect 48190 7520 50000 7576
rect 48129 7518 50000 7520
rect 48129 7515 48195 7518
rect 49200 7488 50000 7518
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 0 6898 800 6928
rect 2773 6898 2839 6901
rect 0 6896 2839 6898
rect 0 6840 2778 6896
rect 2834 6840 2839 6896
rect 0 6838 2839 6840
rect 0 6808 800 6838
rect 2773 6835 2839 6838
rect 45553 6898 45619 6901
rect 49200 6898 50000 6928
rect 45553 6896 50000 6898
rect 45553 6840 45558 6896
rect 45614 6840 50000 6896
rect 45553 6838 50000 6840
rect 45553 6835 45619 6838
rect 49200 6808 50000 6838
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 0 6218 800 6248
rect 3417 6218 3483 6221
rect 0 6216 3483 6218
rect 0 6160 3422 6216
rect 3478 6160 3483 6216
rect 0 6158 3483 6160
rect 0 6128 800 6158
rect 3417 6155 3483 6158
rect 45645 6218 45711 6221
rect 49200 6218 50000 6248
rect 45645 6216 50000 6218
rect 45645 6160 45650 6216
rect 45706 6160 50000 6216
rect 45645 6158 50000 6160
rect 45645 6155 45711 6158
rect 49200 6128 50000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 0 5538 800 5568
rect 2773 5538 2839 5541
rect 0 5536 2839 5538
rect 0 5480 2778 5536
rect 2834 5480 2839 5536
rect 0 5478 2839 5480
rect 0 5448 800 5478
rect 2773 5475 2839 5478
rect 47945 5538 48011 5541
rect 49200 5538 50000 5568
rect 47945 5536 50000 5538
rect 47945 5480 47950 5536
rect 48006 5480 50000 5536
rect 47945 5478 50000 5480
rect 47945 5475 48011 5478
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 49200 5448 50000 5478
rect 19568 5407 19888 5408
rect 4208 4928 4528 4929
rect 0 4858 800 4888
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 3233 4858 3299 4861
rect 0 4856 3299 4858
rect 0 4800 3238 4856
rect 3294 4800 3299 4856
rect 0 4798 3299 4800
rect 0 4768 800 4798
rect 3233 4795 3299 4798
rect 48129 4858 48195 4861
rect 49200 4858 50000 4888
rect 48129 4856 50000 4858
rect 48129 4800 48134 4856
rect 48190 4800 50000 4856
rect 48129 4798 50000 4800
rect 48129 4795 48195 4798
rect 49200 4768 50000 4798
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 0 4178 800 4208
rect 3417 4178 3483 4181
rect 0 4176 3483 4178
rect 0 4120 3422 4176
rect 3478 4120 3483 4176
rect 0 4118 3483 4120
rect 0 4088 800 4118
rect 3417 4115 3483 4118
rect 46197 4178 46263 4181
rect 49200 4178 50000 4208
rect 46197 4176 50000 4178
rect 46197 4120 46202 4176
rect 46258 4120 50000 4176
rect 46197 4118 50000 4120
rect 46197 4115 46263 4118
rect 49200 4088 50000 4118
rect 12433 4042 12499 4045
rect 17677 4042 17743 4045
rect 12433 4040 17743 4042
rect 12433 3984 12438 4040
rect 12494 3984 17682 4040
rect 17738 3984 17743 4040
rect 12433 3982 17743 3984
rect 12433 3979 12499 3982
rect 17677 3979 17743 3982
rect 22553 4042 22619 4045
rect 24393 4042 24459 4045
rect 22553 4040 24459 4042
rect 22553 3984 22558 4040
rect 22614 3984 24398 4040
rect 24454 3984 24459 4040
rect 22553 3982 24459 3984
rect 22553 3979 22619 3982
rect 24393 3979 24459 3982
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 0 3498 800 3528
rect 1853 3498 1919 3501
rect 0 3496 1919 3498
rect 0 3440 1858 3496
rect 1914 3440 1919 3496
rect 0 3438 1919 3440
rect 0 3408 800 3438
rect 1853 3435 1919 3438
rect 45553 3498 45619 3501
rect 49200 3498 50000 3528
rect 45553 3496 50000 3498
rect 45553 3440 45558 3496
rect 45614 3440 50000 3496
rect 45553 3438 50000 3440
rect 45553 3435 45619 3438
rect 49200 3408 50000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 30189 2954 30255 2957
rect 31293 2954 31359 2957
rect 30189 2952 31359 2954
rect 30189 2896 30194 2952
rect 30250 2896 31298 2952
rect 31354 2896 31359 2952
rect 30189 2894 31359 2896
rect 30189 2891 30255 2894
rect 31293 2891 31359 2894
rect 0 2728 800 2848
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 49200 2728 50000 2848
rect 34928 2687 35248 2688
rect 23974 2484 23980 2548
rect 24044 2546 24050 2548
rect 35065 2546 35131 2549
rect 24044 2544 35131 2546
rect 24044 2488 35070 2544
rect 35126 2488 35131 2544
rect 24044 2486 35131 2488
rect 24044 2484 24050 2486
rect 35065 2483 35131 2486
rect 4797 2410 4863 2413
rect 24526 2410 24532 2412
rect 4797 2408 24532 2410
rect 4797 2352 4802 2408
rect 4858 2352 24532 2408
rect 4797 2350 24532 2352
rect 4797 2347 4863 2350
rect 24526 2348 24532 2350
rect 24596 2348 24602 2412
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 4061 2138 4127 2141
rect 0 2136 4127 2138
rect 0 2080 4066 2136
rect 4122 2080 4127 2136
rect 0 2078 4127 2080
rect 0 2048 800 2078
rect 4061 2075 4127 2078
rect 49200 2048 50000 2168
rect 0 1368 800 1488
rect 46841 1458 46907 1461
rect 49200 1458 50000 1488
rect 46841 1456 50000 1458
rect 46841 1400 46846 1456
rect 46902 1400 50000 1456
rect 46841 1398 50000 1400
rect 46841 1395 46907 1398
rect 49200 1368 50000 1398
rect 0 778 800 808
rect 2773 778 2839 781
rect 0 776 2839 778
rect 0 720 2778 776
rect 2834 720 2839 776
rect 0 718 2839 720
rect 0 688 800 718
rect 2773 715 2839 718
rect 47761 778 47827 781
rect 49200 778 50000 808
rect 47761 776 50000 778
rect 47761 720 47766 776
rect 47822 720 50000 776
rect 47761 718 50000 720
rect 47761 715 47827 718
rect 49200 688 50000 718
rect 46749 98 46815 101
rect 49200 98 50000 128
rect 46749 96 50000 98
rect 46749 40 46754 96
rect 46810 40 50000 96
rect 46749 38 50000 40
rect 46749 35 46815 38
rect 49200 8 50000 38
<< via3 >>
rect 4216 49532 4280 49536
rect 4216 49476 4220 49532
rect 4220 49476 4276 49532
rect 4276 49476 4280 49532
rect 4216 49472 4280 49476
rect 4296 49532 4360 49536
rect 4296 49476 4300 49532
rect 4300 49476 4356 49532
rect 4356 49476 4360 49532
rect 4296 49472 4360 49476
rect 4376 49532 4440 49536
rect 4376 49476 4380 49532
rect 4380 49476 4436 49532
rect 4436 49476 4440 49532
rect 4376 49472 4440 49476
rect 4456 49532 4520 49536
rect 4456 49476 4460 49532
rect 4460 49476 4516 49532
rect 4516 49476 4520 49532
rect 4456 49472 4520 49476
rect 34936 49532 35000 49536
rect 34936 49476 34940 49532
rect 34940 49476 34996 49532
rect 34996 49476 35000 49532
rect 34936 49472 35000 49476
rect 35016 49532 35080 49536
rect 35016 49476 35020 49532
rect 35020 49476 35076 49532
rect 35076 49476 35080 49532
rect 35016 49472 35080 49476
rect 35096 49532 35160 49536
rect 35096 49476 35100 49532
rect 35100 49476 35156 49532
rect 35156 49476 35160 49532
rect 35096 49472 35160 49476
rect 35176 49532 35240 49536
rect 35176 49476 35180 49532
rect 35180 49476 35236 49532
rect 35236 49476 35240 49532
rect 35176 49472 35240 49476
rect 19576 48988 19640 48992
rect 19576 48932 19580 48988
rect 19580 48932 19636 48988
rect 19636 48932 19640 48988
rect 19576 48928 19640 48932
rect 19656 48988 19720 48992
rect 19656 48932 19660 48988
rect 19660 48932 19716 48988
rect 19716 48932 19720 48988
rect 19656 48928 19720 48932
rect 19736 48988 19800 48992
rect 19736 48932 19740 48988
rect 19740 48932 19796 48988
rect 19796 48932 19800 48988
rect 19736 48928 19800 48932
rect 19816 48988 19880 48992
rect 19816 48932 19820 48988
rect 19820 48932 19876 48988
rect 19876 48932 19880 48988
rect 19816 48928 19880 48932
rect 4216 48444 4280 48448
rect 4216 48388 4220 48444
rect 4220 48388 4276 48444
rect 4276 48388 4280 48444
rect 4216 48384 4280 48388
rect 4296 48444 4360 48448
rect 4296 48388 4300 48444
rect 4300 48388 4356 48444
rect 4356 48388 4360 48444
rect 4296 48384 4360 48388
rect 4376 48444 4440 48448
rect 4376 48388 4380 48444
rect 4380 48388 4436 48444
rect 4436 48388 4440 48444
rect 4376 48384 4440 48388
rect 4456 48444 4520 48448
rect 4456 48388 4460 48444
rect 4460 48388 4516 48444
rect 4516 48388 4520 48444
rect 4456 48384 4520 48388
rect 34936 48444 35000 48448
rect 34936 48388 34940 48444
rect 34940 48388 34996 48444
rect 34996 48388 35000 48444
rect 34936 48384 35000 48388
rect 35016 48444 35080 48448
rect 35016 48388 35020 48444
rect 35020 48388 35076 48444
rect 35076 48388 35080 48444
rect 35016 48384 35080 48388
rect 35096 48444 35160 48448
rect 35096 48388 35100 48444
rect 35100 48388 35156 48444
rect 35156 48388 35160 48444
rect 35096 48384 35160 48388
rect 35176 48444 35240 48448
rect 35176 48388 35180 48444
rect 35180 48388 35236 48444
rect 35236 48388 35240 48444
rect 35176 48384 35240 48388
rect 19576 47900 19640 47904
rect 19576 47844 19580 47900
rect 19580 47844 19636 47900
rect 19636 47844 19640 47900
rect 19576 47840 19640 47844
rect 19656 47900 19720 47904
rect 19656 47844 19660 47900
rect 19660 47844 19716 47900
rect 19716 47844 19720 47900
rect 19656 47840 19720 47844
rect 19736 47900 19800 47904
rect 19736 47844 19740 47900
rect 19740 47844 19796 47900
rect 19796 47844 19800 47900
rect 19736 47840 19800 47844
rect 19816 47900 19880 47904
rect 19816 47844 19820 47900
rect 19820 47844 19876 47900
rect 19876 47844 19880 47900
rect 19816 47840 19880 47844
rect 4216 47356 4280 47360
rect 4216 47300 4220 47356
rect 4220 47300 4276 47356
rect 4276 47300 4280 47356
rect 4216 47296 4280 47300
rect 4296 47356 4360 47360
rect 4296 47300 4300 47356
rect 4300 47300 4356 47356
rect 4356 47300 4360 47356
rect 4296 47296 4360 47300
rect 4376 47356 4440 47360
rect 4376 47300 4380 47356
rect 4380 47300 4436 47356
rect 4436 47300 4440 47356
rect 4376 47296 4440 47300
rect 4456 47356 4520 47360
rect 4456 47300 4460 47356
rect 4460 47300 4516 47356
rect 4516 47300 4520 47356
rect 4456 47296 4520 47300
rect 34936 47356 35000 47360
rect 34936 47300 34940 47356
rect 34940 47300 34996 47356
rect 34996 47300 35000 47356
rect 34936 47296 35000 47300
rect 35016 47356 35080 47360
rect 35016 47300 35020 47356
rect 35020 47300 35076 47356
rect 35076 47300 35080 47356
rect 35016 47296 35080 47300
rect 35096 47356 35160 47360
rect 35096 47300 35100 47356
rect 35100 47300 35156 47356
rect 35156 47300 35160 47356
rect 35096 47296 35160 47300
rect 35176 47356 35240 47360
rect 35176 47300 35180 47356
rect 35180 47300 35236 47356
rect 35236 47300 35240 47356
rect 35176 47296 35240 47300
rect 19576 46812 19640 46816
rect 19576 46756 19580 46812
rect 19580 46756 19636 46812
rect 19636 46756 19640 46812
rect 19576 46752 19640 46756
rect 19656 46812 19720 46816
rect 19656 46756 19660 46812
rect 19660 46756 19716 46812
rect 19716 46756 19720 46812
rect 19656 46752 19720 46756
rect 19736 46812 19800 46816
rect 19736 46756 19740 46812
rect 19740 46756 19796 46812
rect 19796 46756 19800 46812
rect 19736 46752 19800 46756
rect 19816 46812 19880 46816
rect 19816 46756 19820 46812
rect 19820 46756 19876 46812
rect 19876 46756 19880 46812
rect 19816 46752 19880 46756
rect 4216 46268 4280 46272
rect 4216 46212 4220 46268
rect 4220 46212 4276 46268
rect 4276 46212 4280 46268
rect 4216 46208 4280 46212
rect 4296 46268 4360 46272
rect 4296 46212 4300 46268
rect 4300 46212 4356 46268
rect 4356 46212 4360 46268
rect 4296 46208 4360 46212
rect 4376 46268 4440 46272
rect 4376 46212 4380 46268
rect 4380 46212 4436 46268
rect 4436 46212 4440 46268
rect 4376 46208 4440 46212
rect 4456 46268 4520 46272
rect 4456 46212 4460 46268
rect 4460 46212 4516 46268
rect 4516 46212 4520 46268
rect 4456 46208 4520 46212
rect 34936 46268 35000 46272
rect 34936 46212 34940 46268
rect 34940 46212 34996 46268
rect 34996 46212 35000 46268
rect 34936 46208 35000 46212
rect 35016 46268 35080 46272
rect 35016 46212 35020 46268
rect 35020 46212 35076 46268
rect 35076 46212 35080 46268
rect 35016 46208 35080 46212
rect 35096 46268 35160 46272
rect 35096 46212 35100 46268
rect 35100 46212 35156 46268
rect 35156 46212 35160 46268
rect 35096 46208 35160 46212
rect 35176 46268 35240 46272
rect 35176 46212 35180 46268
rect 35180 46212 35236 46268
rect 35236 46212 35240 46268
rect 35176 46208 35240 46212
rect 19576 45724 19640 45728
rect 19576 45668 19580 45724
rect 19580 45668 19636 45724
rect 19636 45668 19640 45724
rect 19576 45664 19640 45668
rect 19656 45724 19720 45728
rect 19656 45668 19660 45724
rect 19660 45668 19716 45724
rect 19716 45668 19720 45724
rect 19656 45664 19720 45668
rect 19736 45724 19800 45728
rect 19736 45668 19740 45724
rect 19740 45668 19796 45724
rect 19796 45668 19800 45724
rect 19736 45664 19800 45668
rect 19816 45724 19880 45728
rect 19816 45668 19820 45724
rect 19820 45668 19876 45724
rect 19876 45668 19880 45724
rect 19816 45664 19880 45668
rect 4216 45180 4280 45184
rect 4216 45124 4220 45180
rect 4220 45124 4276 45180
rect 4276 45124 4280 45180
rect 4216 45120 4280 45124
rect 4296 45180 4360 45184
rect 4296 45124 4300 45180
rect 4300 45124 4356 45180
rect 4356 45124 4360 45180
rect 4296 45120 4360 45124
rect 4376 45180 4440 45184
rect 4376 45124 4380 45180
rect 4380 45124 4436 45180
rect 4436 45124 4440 45180
rect 4376 45120 4440 45124
rect 4456 45180 4520 45184
rect 4456 45124 4460 45180
rect 4460 45124 4516 45180
rect 4516 45124 4520 45180
rect 4456 45120 4520 45124
rect 34936 45180 35000 45184
rect 34936 45124 34940 45180
rect 34940 45124 34996 45180
rect 34996 45124 35000 45180
rect 34936 45120 35000 45124
rect 35016 45180 35080 45184
rect 35016 45124 35020 45180
rect 35020 45124 35076 45180
rect 35076 45124 35080 45180
rect 35016 45120 35080 45124
rect 35096 45180 35160 45184
rect 35096 45124 35100 45180
rect 35100 45124 35156 45180
rect 35156 45124 35160 45180
rect 35096 45120 35160 45124
rect 35176 45180 35240 45184
rect 35176 45124 35180 45180
rect 35180 45124 35236 45180
rect 35236 45124 35240 45180
rect 35176 45120 35240 45124
rect 19576 44636 19640 44640
rect 19576 44580 19580 44636
rect 19580 44580 19636 44636
rect 19636 44580 19640 44636
rect 19576 44576 19640 44580
rect 19656 44636 19720 44640
rect 19656 44580 19660 44636
rect 19660 44580 19716 44636
rect 19716 44580 19720 44636
rect 19656 44576 19720 44580
rect 19736 44636 19800 44640
rect 19736 44580 19740 44636
rect 19740 44580 19796 44636
rect 19796 44580 19800 44636
rect 19736 44576 19800 44580
rect 19816 44636 19880 44640
rect 19816 44580 19820 44636
rect 19820 44580 19876 44636
rect 19876 44580 19880 44636
rect 19816 44576 19880 44580
rect 4216 44092 4280 44096
rect 4216 44036 4220 44092
rect 4220 44036 4276 44092
rect 4276 44036 4280 44092
rect 4216 44032 4280 44036
rect 4296 44092 4360 44096
rect 4296 44036 4300 44092
rect 4300 44036 4356 44092
rect 4356 44036 4360 44092
rect 4296 44032 4360 44036
rect 4376 44092 4440 44096
rect 4376 44036 4380 44092
rect 4380 44036 4436 44092
rect 4436 44036 4440 44092
rect 4376 44032 4440 44036
rect 4456 44092 4520 44096
rect 4456 44036 4460 44092
rect 4460 44036 4516 44092
rect 4516 44036 4520 44092
rect 4456 44032 4520 44036
rect 34936 44092 35000 44096
rect 34936 44036 34940 44092
rect 34940 44036 34996 44092
rect 34996 44036 35000 44092
rect 34936 44032 35000 44036
rect 35016 44092 35080 44096
rect 35016 44036 35020 44092
rect 35020 44036 35076 44092
rect 35076 44036 35080 44092
rect 35016 44032 35080 44036
rect 35096 44092 35160 44096
rect 35096 44036 35100 44092
rect 35100 44036 35156 44092
rect 35156 44036 35160 44092
rect 35096 44032 35160 44036
rect 35176 44092 35240 44096
rect 35176 44036 35180 44092
rect 35180 44036 35236 44092
rect 35236 44036 35240 44092
rect 35176 44032 35240 44036
rect 19576 43548 19640 43552
rect 19576 43492 19580 43548
rect 19580 43492 19636 43548
rect 19636 43492 19640 43548
rect 19576 43488 19640 43492
rect 19656 43548 19720 43552
rect 19656 43492 19660 43548
rect 19660 43492 19716 43548
rect 19716 43492 19720 43548
rect 19656 43488 19720 43492
rect 19736 43548 19800 43552
rect 19736 43492 19740 43548
rect 19740 43492 19796 43548
rect 19796 43492 19800 43548
rect 19736 43488 19800 43492
rect 19816 43548 19880 43552
rect 19816 43492 19820 43548
rect 19820 43492 19876 43548
rect 19876 43492 19880 43548
rect 19816 43488 19880 43492
rect 4216 43004 4280 43008
rect 4216 42948 4220 43004
rect 4220 42948 4276 43004
rect 4276 42948 4280 43004
rect 4216 42944 4280 42948
rect 4296 43004 4360 43008
rect 4296 42948 4300 43004
rect 4300 42948 4356 43004
rect 4356 42948 4360 43004
rect 4296 42944 4360 42948
rect 4376 43004 4440 43008
rect 4376 42948 4380 43004
rect 4380 42948 4436 43004
rect 4436 42948 4440 43004
rect 4376 42944 4440 42948
rect 4456 43004 4520 43008
rect 4456 42948 4460 43004
rect 4460 42948 4516 43004
rect 4516 42948 4520 43004
rect 4456 42944 4520 42948
rect 34936 43004 35000 43008
rect 34936 42948 34940 43004
rect 34940 42948 34996 43004
rect 34996 42948 35000 43004
rect 34936 42944 35000 42948
rect 35016 43004 35080 43008
rect 35016 42948 35020 43004
rect 35020 42948 35076 43004
rect 35076 42948 35080 43004
rect 35016 42944 35080 42948
rect 35096 43004 35160 43008
rect 35096 42948 35100 43004
rect 35100 42948 35156 43004
rect 35156 42948 35160 43004
rect 35096 42944 35160 42948
rect 35176 43004 35240 43008
rect 35176 42948 35180 43004
rect 35180 42948 35236 43004
rect 35236 42948 35240 43004
rect 35176 42944 35240 42948
rect 19576 42460 19640 42464
rect 19576 42404 19580 42460
rect 19580 42404 19636 42460
rect 19636 42404 19640 42460
rect 19576 42400 19640 42404
rect 19656 42460 19720 42464
rect 19656 42404 19660 42460
rect 19660 42404 19716 42460
rect 19716 42404 19720 42460
rect 19656 42400 19720 42404
rect 19736 42460 19800 42464
rect 19736 42404 19740 42460
rect 19740 42404 19796 42460
rect 19796 42404 19800 42460
rect 19736 42400 19800 42404
rect 19816 42460 19880 42464
rect 19816 42404 19820 42460
rect 19820 42404 19876 42460
rect 19876 42404 19880 42460
rect 19816 42400 19880 42404
rect 4216 41916 4280 41920
rect 4216 41860 4220 41916
rect 4220 41860 4276 41916
rect 4276 41860 4280 41916
rect 4216 41856 4280 41860
rect 4296 41916 4360 41920
rect 4296 41860 4300 41916
rect 4300 41860 4356 41916
rect 4356 41860 4360 41916
rect 4296 41856 4360 41860
rect 4376 41916 4440 41920
rect 4376 41860 4380 41916
rect 4380 41860 4436 41916
rect 4436 41860 4440 41916
rect 4376 41856 4440 41860
rect 4456 41916 4520 41920
rect 4456 41860 4460 41916
rect 4460 41860 4516 41916
rect 4516 41860 4520 41916
rect 4456 41856 4520 41860
rect 34936 41916 35000 41920
rect 34936 41860 34940 41916
rect 34940 41860 34996 41916
rect 34996 41860 35000 41916
rect 34936 41856 35000 41860
rect 35016 41916 35080 41920
rect 35016 41860 35020 41916
rect 35020 41860 35076 41916
rect 35076 41860 35080 41916
rect 35016 41856 35080 41860
rect 35096 41916 35160 41920
rect 35096 41860 35100 41916
rect 35100 41860 35156 41916
rect 35156 41860 35160 41916
rect 35096 41856 35160 41860
rect 35176 41916 35240 41920
rect 35176 41860 35180 41916
rect 35180 41860 35236 41916
rect 35236 41860 35240 41916
rect 35176 41856 35240 41860
rect 19576 41372 19640 41376
rect 19576 41316 19580 41372
rect 19580 41316 19636 41372
rect 19636 41316 19640 41372
rect 19576 41312 19640 41316
rect 19656 41372 19720 41376
rect 19656 41316 19660 41372
rect 19660 41316 19716 41372
rect 19716 41316 19720 41372
rect 19656 41312 19720 41316
rect 19736 41372 19800 41376
rect 19736 41316 19740 41372
rect 19740 41316 19796 41372
rect 19796 41316 19800 41372
rect 19736 41312 19800 41316
rect 19816 41372 19880 41376
rect 19816 41316 19820 41372
rect 19820 41316 19876 41372
rect 19876 41316 19880 41372
rect 19816 41312 19880 41316
rect 4216 40828 4280 40832
rect 4216 40772 4220 40828
rect 4220 40772 4276 40828
rect 4276 40772 4280 40828
rect 4216 40768 4280 40772
rect 4296 40828 4360 40832
rect 4296 40772 4300 40828
rect 4300 40772 4356 40828
rect 4356 40772 4360 40828
rect 4296 40768 4360 40772
rect 4376 40828 4440 40832
rect 4376 40772 4380 40828
rect 4380 40772 4436 40828
rect 4436 40772 4440 40828
rect 4376 40768 4440 40772
rect 4456 40828 4520 40832
rect 4456 40772 4460 40828
rect 4460 40772 4516 40828
rect 4516 40772 4520 40828
rect 4456 40768 4520 40772
rect 34936 40828 35000 40832
rect 34936 40772 34940 40828
rect 34940 40772 34996 40828
rect 34996 40772 35000 40828
rect 34936 40768 35000 40772
rect 35016 40828 35080 40832
rect 35016 40772 35020 40828
rect 35020 40772 35076 40828
rect 35076 40772 35080 40828
rect 35016 40768 35080 40772
rect 35096 40828 35160 40832
rect 35096 40772 35100 40828
rect 35100 40772 35156 40828
rect 35156 40772 35160 40828
rect 35096 40768 35160 40772
rect 35176 40828 35240 40832
rect 35176 40772 35180 40828
rect 35180 40772 35236 40828
rect 35236 40772 35240 40828
rect 35176 40768 35240 40772
rect 19576 40284 19640 40288
rect 19576 40228 19580 40284
rect 19580 40228 19636 40284
rect 19636 40228 19640 40284
rect 19576 40224 19640 40228
rect 19656 40284 19720 40288
rect 19656 40228 19660 40284
rect 19660 40228 19716 40284
rect 19716 40228 19720 40284
rect 19656 40224 19720 40228
rect 19736 40284 19800 40288
rect 19736 40228 19740 40284
rect 19740 40228 19796 40284
rect 19796 40228 19800 40284
rect 19736 40224 19800 40228
rect 19816 40284 19880 40288
rect 19816 40228 19820 40284
rect 19820 40228 19876 40284
rect 19876 40228 19880 40284
rect 19816 40224 19880 40228
rect 4216 39740 4280 39744
rect 4216 39684 4220 39740
rect 4220 39684 4276 39740
rect 4276 39684 4280 39740
rect 4216 39680 4280 39684
rect 4296 39740 4360 39744
rect 4296 39684 4300 39740
rect 4300 39684 4356 39740
rect 4356 39684 4360 39740
rect 4296 39680 4360 39684
rect 4376 39740 4440 39744
rect 4376 39684 4380 39740
rect 4380 39684 4436 39740
rect 4436 39684 4440 39740
rect 4376 39680 4440 39684
rect 4456 39740 4520 39744
rect 4456 39684 4460 39740
rect 4460 39684 4516 39740
rect 4516 39684 4520 39740
rect 4456 39680 4520 39684
rect 34936 39740 35000 39744
rect 34936 39684 34940 39740
rect 34940 39684 34996 39740
rect 34996 39684 35000 39740
rect 34936 39680 35000 39684
rect 35016 39740 35080 39744
rect 35016 39684 35020 39740
rect 35020 39684 35076 39740
rect 35076 39684 35080 39740
rect 35016 39680 35080 39684
rect 35096 39740 35160 39744
rect 35096 39684 35100 39740
rect 35100 39684 35156 39740
rect 35156 39684 35160 39740
rect 35096 39680 35160 39684
rect 35176 39740 35240 39744
rect 35176 39684 35180 39740
rect 35180 39684 35236 39740
rect 35236 39684 35240 39740
rect 35176 39680 35240 39684
rect 19576 39196 19640 39200
rect 19576 39140 19580 39196
rect 19580 39140 19636 39196
rect 19636 39140 19640 39196
rect 19576 39136 19640 39140
rect 19656 39196 19720 39200
rect 19656 39140 19660 39196
rect 19660 39140 19716 39196
rect 19716 39140 19720 39196
rect 19656 39136 19720 39140
rect 19736 39196 19800 39200
rect 19736 39140 19740 39196
rect 19740 39140 19796 39196
rect 19796 39140 19800 39196
rect 19736 39136 19800 39140
rect 19816 39196 19880 39200
rect 19816 39140 19820 39196
rect 19820 39140 19876 39196
rect 19876 39140 19880 39196
rect 19816 39136 19880 39140
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 19576 38108 19640 38112
rect 19576 38052 19580 38108
rect 19580 38052 19636 38108
rect 19636 38052 19640 38108
rect 19576 38048 19640 38052
rect 19656 38108 19720 38112
rect 19656 38052 19660 38108
rect 19660 38052 19716 38108
rect 19716 38052 19720 38108
rect 19656 38048 19720 38052
rect 19736 38108 19800 38112
rect 19736 38052 19740 38108
rect 19740 38052 19796 38108
rect 19796 38052 19800 38108
rect 19736 38048 19800 38052
rect 19816 38108 19880 38112
rect 19816 38052 19820 38108
rect 19820 38052 19876 38108
rect 19876 38052 19880 38108
rect 19816 38048 19880 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 20116 33008 20180 33012
rect 20116 32952 20166 33008
rect 20166 32952 20180 33008
rect 20116 32948 20180 32952
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 23428 30228 23492 30292
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 20116 29140 20180 29204
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 24348 25060 24412 25124
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 23428 22884 23492 22948
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 24532 20708 24596 20772
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 24348 20436 24412 20500
rect 23980 20300 24044 20364
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 28212 17776 28276 17780
rect 28212 17720 28226 17776
rect 28226 17720 28276 17776
rect 28212 17716 28276 17720
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 28212 16356 28276 16420
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 23980 2484 24044 2548
rect 24532 2348 24596 2412
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
<< metal4 >>
rect 4208 49536 4528 49552
rect 4208 49472 4216 49536
rect 4280 49472 4296 49536
rect 4360 49472 4376 49536
rect 4440 49472 4456 49536
rect 4520 49472 4528 49536
rect 4208 48448 4528 49472
rect 4208 48384 4216 48448
rect 4280 48384 4296 48448
rect 4360 48384 4376 48448
rect 4440 48384 4456 48448
rect 4520 48384 4528 48448
rect 4208 47360 4528 48384
rect 4208 47296 4216 47360
rect 4280 47296 4296 47360
rect 4360 47296 4376 47360
rect 4440 47296 4456 47360
rect 4520 47296 4528 47360
rect 4208 46272 4528 47296
rect 4208 46208 4216 46272
rect 4280 46208 4296 46272
rect 4360 46208 4376 46272
rect 4440 46208 4456 46272
rect 4520 46208 4528 46272
rect 4208 45184 4528 46208
rect 4208 45120 4216 45184
rect 4280 45120 4296 45184
rect 4360 45120 4376 45184
rect 4440 45120 4456 45184
rect 4520 45120 4528 45184
rect 4208 44096 4528 45120
rect 4208 44032 4216 44096
rect 4280 44032 4296 44096
rect 4360 44032 4376 44096
rect 4440 44032 4456 44096
rect 4520 44032 4528 44096
rect 4208 43008 4528 44032
rect 4208 42944 4216 43008
rect 4280 42944 4296 43008
rect 4360 42944 4376 43008
rect 4440 42944 4456 43008
rect 4520 42944 4528 43008
rect 4208 41920 4528 42944
rect 4208 41856 4216 41920
rect 4280 41856 4296 41920
rect 4360 41856 4376 41920
rect 4440 41856 4456 41920
rect 4520 41856 4528 41920
rect 4208 40832 4528 41856
rect 4208 40768 4216 40832
rect 4280 40768 4296 40832
rect 4360 40768 4376 40832
rect 4440 40768 4456 40832
rect 4520 40768 4528 40832
rect 4208 39744 4528 40768
rect 4208 39680 4216 39744
rect 4280 39680 4296 39744
rect 4360 39680 4376 39744
rect 4440 39680 4456 39744
rect 4520 39680 4528 39744
rect 4208 38656 4528 39680
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 48992 19888 49552
rect 19568 48928 19576 48992
rect 19640 48928 19656 48992
rect 19720 48928 19736 48992
rect 19800 48928 19816 48992
rect 19880 48928 19888 48992
rect 19568 47904 19888 48928
rect 19568 47840 19576 47904
rect 19640 47840 19656 47904
rect 19720 47840 19736 47904
rect 19800 47840 19816 47904
rect 19880 47840 19888 47904
rect 19568 46816 19888 47840
rect 19568 46752 19576 46816
rect 19640 46752 19656 46816
rect 19720 46752 19736 46816
rect 19800 46752 19816 46816
rect 19880 46752 19888 46816
rect 19568 45728 19888 46752
rect 19568 45664 19576 45728
rect 19640 45664 19656 45728
rect 19720 45664 19736 45728
rect 19800 45664 19816 45728
rect 19880 45664 19888 45728
rect 19568 44640 19888 45664
rect 19568 44576 19576 44640
rect 19640 44576 19656 44640
rect 19720 44576 19736 44640
rect 19800 44576 19816 44640
rect 19880 44576 19888 44640
rect 19568 43552 19888 44576
rect 19568 43488 19576 43552
rect 19640 43488 19656 43552
rect 19720 43488 19736 43552
rect 19800 43488 19816 43552
rect 19880 43488 19888 43552
rect 19568 42464 19888 43488
rect 19568 42400 19576 42464
rect 19640 42400 19656 42464
rect 19720 42400 19736 42464
rect 19800 42400 19816 42464
rect 19880 42400 19888 42464
rect 19568 41376 19888 42400
rect 19568 41312 19576 41376
rect 19640 41312 19656 41376
rect 19720 41312 19736 41376
rect 19800 41312 19816 41376
rect 19880 41312 19888 41376
rect 19568 40288 19888 41312
rect 19568 40224 19576 40288
rect 19640 40224 19656 40288
rect 19720 40224 19736 40288
rect 19800 40224 19816 40288
rect 19880 40224 19888 40288
rect 19568 39200 19888 40224
rect 19568 39136 19576 39200
rect 19640 39136 19656 39200
rect 19720 39136 19736 39200
rect 19800 39136 19816 39200
rect 19880 39136 19888 39200
rect 19568 38112 19888 39136
rect 19568 38048 19576 38112
rect 19640 38048 19656 38112
rect 19720 38048 19736 38112
rect 19800 38048 19816 38112
rect 19880 38048 19888 38112
rect 19568 37024 19888 38048
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 34928 49536 35248 49552
rect 34928 49472 34936 49536
rect 35000 49472 35016 49536
rect 35080 49472 35096 49536
rect 35160 49472 35176 49536
rect 35240 49472 35248 49536
rect 34928 48448 35248 49472
rect 34928 48384 34936 48448
rect 35000 48384 35016 48448
rect 35080 48384 35096 48448
rect 35160 48384 35176 48448
rect 35240 48384 35248 48448
rect 34928 47360 35248 48384
rect 34928 47296 34936 47360
rect 35000 47296 35016 47360
rect 35080 47296 35096 47360
rect 35160 47296 35176 47360
rect 35240 47296 35248 47360
rect 34928 46272 35248 47296
rect 34928 46208 34936 46272
rect 35000 46208 35016 46272
rect 35080 46208 35096 46272
rect 35160 46208 35176 46272
rect 35240 46208 35248 46272
rect 34928 45184 35248 46208
rect 34928 45120 34936 45184
rect 35000 45120 35016 45184
rect 35080 45120 35096 45184
rect 35160 45120 35176 45184
rect 35240 45120 35248 45184
rect 34928 44096 35248 45120
rect 34928 44032 34936 44096
rect 35000 44032 35016 44096
rect 35080 44032 35096 44096
rect 35160 44032 35176 44096
rect 35240 44032 35248 44096
rect 34928 43008 35248 44032
rect 34928 42944 34936 43008
rect 35000 42944 35016 43008
rect 35080 42944 35096 43008
rect 35160 42944 35176 43008
rect 35240 42944 35248 43008
rect 34928 41920 35248 42944
rect 34928 41856 34936 41920
rect 35000 41856 35016 41920
rect 35080 41856 35096 41920
rect 35160 41856 35176 41920
rect 35240 41856 35248 41920
rect 34928 40832 35248 41856
rect 34928 40768 34936 40832
rect 35000 40768 35016 40832
rect 35080 40768 35096 40832
rect 35160 40768 35176 40832
rect 35240 40768 35248 40832
rect 34928 39744 35248 40768
rect 34928 39680 34936 39744
rect 35000 39680 35016 39744
rect 35080 39680 35096 39744
rect 35160 39680 35176 39744
rect 35240 39680 35248 39744
rect 34928 38656 35248 39680
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 20115 33012 20181 33013
rect 20115 32948 20116 33012
rect 20180 32948 20181 33012
rect 20115 32947 20181 32948
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 20118 29205 20178 32947
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 23427 30292 23493 30293
rect 23427 30228 23428 30292
rect 23492 30228 23493 30292
rect 23427 30227 23493 30228
rect 20115 29204 20181 29205
rect 20115 29140 20116 29204
rect 20180 29140 20181 29204
rect 20115 29139 20181 29140
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 23430 22949 23490 30227
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 24347 25124 24413 25125
rect 24347 25060 24348 25124
rect 24412 25060 24413 25124
rect 24347 25059 24413 25060
rect 23427 22948 23493 22949
rect 23427 22884 23428 22948
rect 23492 22884 23493 22948
rect 23427 22883 23493 22884
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 24350 20501 24410 25059
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 24531 20772 24597 20773
rect 24531 20708 24532 20772
rect 24596 20708 24597 20772
rect 24531 20707 24597 20708
rect 24347 20500 24413 20501
rect 24347 20436 24348 20500
rect 24412 20436 24413 20500
rect 24347 20435 24413 20436
rect 23979 20364 24045 20365
rect 23979 20300 23980 20364
rect 24044 20300 24045 20364
rect 23979 20299 24045 20300
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 23982 2549 24042 20299
rect 23979 2548 24045 2549
rect 23979 2484 23980 2548
rect 24044 2484 24045 2548
rect 23979 2483 24045 2484
rect 24534 2413 24594 20707
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 28211 17780 28277 17781
rect 28211 17716 28212 17780
rect 28276 17716 28277 17780
rect 28211 17715 28277 17716
rect 28214 16421 28274 17715
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 28211 16420 28277 16421
rect 28211 16356 28212 16420
rect 28276 16356 28277 16420
rect 28211 16355 28277 16356
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 24531 2412 24597 2413
rect 24531 2348 24532 2412
rect 24596 2348 24597 2412
rect 24531 2347 24597 2348
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 2128 35248 2688
use sky130_fd_sc_hd__diode_2  ANTENNA_0 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 17296 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1
timestamp 1644511149
transform 1 0 41860 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1644511149
transform 1 0 22632 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1644511149
transform 1 0 27784 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1644511149
transform 1 0 7176 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1644511149
transform 1 0 24288 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1644511149
transform 1 0 24656 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1644511149
transform 1 0 17572 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3312 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4048 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_0_42 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4968 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_78
timestamp 1644511149
transform 1 0 8280 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_95
timestamp 1644511149
transform 1 0 9844 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_105
timestamp 1644511149
transform 1 0 10764 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_111 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11316 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_113 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_121 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 12236 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_127
timestamp 1644511149
transform 1 0 12788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_134
timestamp 1644511149
transform 1 0 13432 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_141
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_149
timestamp 1644511149
transform 1 0 14812 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_161
timestamp 1644511149
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_167
timestamp 1644511149
transform 1 0 16468 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_169
timestamp 1644511149
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_177
timestamp 1644511149
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_182
timestamp 1644511149
transform 1 0 17848 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_194
timestamp 1644511149
transform 1 0 18952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_205
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_210
timestamp 1644511149
transform 1 0 20424 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_222
timestamp 1644511149
transform 1 0 21528 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_246
timestamp 1644511149
transform 1 0 23736 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_265
timestamp 1644511149
transform 1 0 25484 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_272
timestamp 1644511149
transform 1 0 26128 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_281
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_286
timestamp 1644511149
transform 1 0 27416 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_300
timestamp 1644511149
transform 1 0 28704 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_345
timestamp 1644511149
transform 1 0 32844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_350
timestamp 1644511149
transform 1 0 33304 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_365
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_371
timestamp 1644511149
transform 1 0 35236 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_379
timestamp 1644511149
transform 1 0 35972 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_384
timestamp 1644511149
transform 1 0 36432 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_405
timestamp 1644511149
transform 1 0 38364 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_416
timestamp 1644511149
transform 1 0 39376 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_433
timestamp 1644511149
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_445
timestamp 1644511149
transform 1 0 42044 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_449
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_457
timestamp 1644511149
transform 1 0 43148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_462
timestamp 1644511149
transform 1 0 43608 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_472
timestamp 1644511149
transform 1 0 44528 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_500
timestamp 1644511149
transform 1 0 47104 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_512
timestamp 1644511149
transform 1 0 48208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_11
timestamp 1644511149
transform 1 0 2116 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_19
timestamp 1644511149
transform 1 0 2852 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_25
timestamp 1644511149
transform 1 0 3404 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_47
timestamp 1644511149
transform 1 0 5428 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_55
timestamp 1644511149
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_78
timestamp 1644511149
transform 1 0 8280 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_92
timestamp 1644511149
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_100
timestamp 1644511149
transform 1 0 10304 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_1_113
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_119
timestamp 1644511149
transform 1 0 12052 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_144
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_1_155
timestamp 1644511149
transform 1 0 15364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_167
timestamp 1644511149
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_169
timestamp 1644511149
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_175
timestamp 1644511149
transform 1 0 17204 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_197
timestamp 1644511149
transform 1 0 19228 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_205
timestamp 1644511149
transform 1 0 19964 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_1_211
timestamp 1644511149
transform 1 0 20516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_1_223
timestamp 1644511149
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_225
timestamp 1644511149
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_233
timestamp 1644511149
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_238
timestamp 1644511149
transform 1 0 23000 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_263
timestamp 1644511149
transform 1 0 25300 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_1_274
timestamp 1644511149
transform 1 0 26312 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_281
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_293
timestamp 1644511149
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_305
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_332
timestamp 1644511149
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_358
timestamp 1644511149
transform 1 0 34040 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_370
timestamp 1644511149
transform 1 0 35144 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_1_378
timestamp 1644511149
transform 1 0 35880 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_383
timestamp 1644511149
transform 1 0 36340 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_391
timestamp 1644511149
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_393
timestamp 1644511149
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_405
timestamp 1644511149
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_1_428
timestamp 1644511149
transform 1 0 40480 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_436
timestamp 1644511149
transform 1 0 41216 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_442
timestamp 1644511149
transform 1 0 41768 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_470
timestamp 1644511149
transform 1 0 44344 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_495
timestamp 1644511149
transform 1 0 46644 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_1_512
timestamp 1644511149
transform 1 0 48208 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_24
timestamp 1644511149
transform 1 0 3312 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_38
timestamp 1644511149
transform 1 0 4600 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_72
timestamp 1644511149
transform 1 0 7728 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_97
timestamp 1644511149
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_109
timestamp 1644511149
transform 1 0 11132 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_136
timestamp 1644511149
transform 1 0 13616 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_141
timestamp 1644511149
transform 1 0 14076 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_148
timestamp 1644511149
transform 1 0 14720 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_173
timestamp 1644511149
transform 1 0 17020 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_179
timestamp 1644511149
transform 1 0 17572 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_183
timestamp 1644511149
transform 1 0 17940 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_2_195
timestamp 1644511149
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_197
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_204
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_229
timestamp 1644511149
transform 1 0 22172 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_233
timestamp 1644511149
transform 1 0 22540 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_237
timestamp 1644511149
transform 1 0 22908 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_244
timestamp 1644511149
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_253
timestamp 1644511149
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_265
timestamp 1644511149
transform 1 0 25484 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_288
timestamp 1644511149
transform 1 0 27600 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_300
timestamp 1644511149
transform 1 0 28704 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_312
timestamp 1644511149
transform 1 0 29808 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_319
timestamp 1644511149
transform 1 0 30452 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_344
timestamp 1644511149
transform 1 0 32752 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_356
timestamp 1644511149
transform 1 0 33856 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_2_401
timestamp 1644511149
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1644511149
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1644511149
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_425
timestamp 1644511149
transform 1 0 40204 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_450
timestamp 1644511149
transform 1 0 42504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_457
timestamp 1644511149
transform 1 0 43148 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_461
timestamp 1644511149
transform 1 0 43516 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_465
timestamp 1644511149
transform 1 0 43884 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_472
timestamp 1644511149
transform 1 0 44528 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_480
timestamp 1644511149
transform 1 0 45264 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_2_509
timestamp 1644511149
transform 1 0 47932 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_515
timestamp 1644511149
transform 1 0 48484 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_6
timestamp 1644511149
transform 1 0 1656 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_13
timestamp 1644511149
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_20
timestamp 1644511149
transform 1 0 2944 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_26
timestamp 1644511149
transform 1 0 3496 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_30
timestamp 1644511149
transform 1 0 3864 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_42
timestamp 1644511149
transform 1 0 4968 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_48
timestamp 1644511149
transform 1 0 5520 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_60
timestamp 1644511149
transform 1 0 6624 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_3_67
timestamp 1644511149
transform 1 0 7268 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_73
timestamp 1644511149
transform 1 0 7820 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_95
timestamp 1644511149
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_107
timestamp 1644511149
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_117
timestamp 1644511149
transform 1 0 11868 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_123
timestamp 1644511149
transform 1 0 12420 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_127
timestamp 1644511149
transform 1 0 12788 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_152
timestamp 1644511149
transform 1 0 15088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_169
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_180
timestamp 1644511149
transform 1 0 17664 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_192
timestamp 1644511149
transform 1 0 18768 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_204
timestamp 1644511149
transform 1 0 19872 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_212
timestamp 1644511149
transform 1 0 20608 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_3_217
timestamp 1644511149
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_223
timestamp 1644511149
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_3_236
timestamp 1644511149
transform 1 0 22816 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_242
timestamp 1644511149
transform 1 0 23368 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_246
timestamp 1644511149
transform 1 0 23736 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_258
timestamp 1644511149
transform 1 0 24840 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_266
timestamp 1644511149
transform 1 0 25576 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_3_271
timestamp 1644511149
transform 1 0 26036 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_279
timestamp 1644511149
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_311
timestamp 1644511149
transform 1 0 29716 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_315
timestamp 1644511149
transform 1 0 30084 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_321
timestamp 1644511149
transform 1 0 30636 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_325
timestamp 1644511149
transform 1 0 31004 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_332
timestamp 1644511149
transform 1 0 31648 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_341
timestamp 1644511149
transform 1 0 32476 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_353
timestamp 1644511149
transform 1 0 33580 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_365
timestamp 1644511149
transform 1 0 34684 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_377
timestamp 1644511149
transform 1 0 35788 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_386
timestamp 1644511149
transform 1 0 36616 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_3_393
timestamp 1644511149
transform 1 0 37260 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_402
timestamp 1644511149
transform 1 0 38088 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_414
timestamp 1644511149
transform 1 0 39192 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_426
timestamp 1644511149
transform 1 0 40296 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_432
timestamp 1644511149
transform 1 0 40848 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_436
timestamp 1644511149
transform 1 0 41216 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_443
timestamp 1644511149
transform 1 0 41860 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_447
timestamp 1644511149
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_452
timestamp 1644511149
transform 1 0 42688 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_3_463
timestamp 1644511149
transform 1 0 43700 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_488
timestamp 1644511149
transform 1 0 46000 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_495
timestamp 1644511149
transform 1 0 46644 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_503
timestamp 1644511149
transform 1 0 47380 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_512
timestamp 1644511149
transform 1 0 48208 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_24
timestamp 1644511149
transform 1 0 3312 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_44
timestamp 1644511149
transform 1 0 5152 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_52
timestamp 1644511149
transform 1 0 5888 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_57
timestamp 1644511149
transform 1 0 6348 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_4_64
timestamp 1644511149
transform 1 0 6992 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_72
timestamp 1644511149
transform 1 0 7728 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_4_78
timestamp 1644511149
transform 1 0 8280 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_97
timestamp 1644511149
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_109
timestamp 1644511149
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_121
timestamp 1644511149
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_133
timestamp 1644511149
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_209
timestamp 1644511149
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_221
timestamp 1644511149
transform 1 0 21436 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_4_248
timestamp 1644511149
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_253
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_265
timestamp 1644511149
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_277
timestamp 1644511149
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_289
timestamp 1644511149
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_301
timestamp 1644511149
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_307
timestamp 1644511149
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_320
timestamp 1644511149
transform 1 0 30544 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_327
timestamp 1644511149
transform 1 0 31188 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_339
timestamp 1644511149
transform 1 0 32292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_351
timestamp 1644511149
transform 1 0 33396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_389
timestamp 1644511149
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_401
timestamp 1644511149
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_413
timestamp 1644511149
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_419
timestamp 1644511149
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_433
timestamp 1644511149
transform 1 0 40940 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_441
timestamp 1644511149
transform 1 0 41676 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_464
timestamp 1644511149
transform 1 0 43792 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_480
timestamp 1644511149
transform 1 0 45264 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_487
timestamp 1644511149
transform 1 0 45908 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_512
timestamp 1644511149
transform 1 0 48208 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_7
timestamp 1644511149
transform 1 0 1748 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_32
timestamp 1644511149
transform 1 0 4048 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_44
timestamp 1644511149
transform 1 0 5152 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_57
timestamp 1644511149
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_69
timestamp 1644511149
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_81
timestamp 1644511149
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_93
timestamp 1644511149
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_105
timestamp 1644511149
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_111
timestamp 1644511149
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_169
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_181
timestamp 1644511149
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_193
timestamp 1644511149
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_205
timestamp 1644511149
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_217
timestamp 1644511149
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_237
timestamp 1644511149
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_249
timestamp 1644511149
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_261
timestamp 1644511149
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_273
timestamp 1644511149
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_279
timestamp 1644511149
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_293
timestamp 1644511149
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_305
timestamp 1644511149
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_317
timestamp 1644511149
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_329
timestamp 1644511149
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_335
timestamp 1644511149
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_349
timestamp 1644511149
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_361
timestamp 1644511149
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_373
timestamp 1644511149
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_385
timestamp 1644511149
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_391
timestamp 1644511149
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_441
timestamp 1644511149
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_447
timestamp 1644511149
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_485
timestamp 1644511149
transform 1 0 45724 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_500
timestamp 1644511149
transform 1 0 47104 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_508
timestamp 1644511149
transform 1 0 47840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_6_14
timestamp 1644511149
transform 1 0 2392 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_6_23
timestamp 1644511149
transform 1 0 3220 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_41
timestamp 1644511149
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_53
timestamp 1644511149
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_65
timestamp 1644511149
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_77
timestamp 1644511149
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_97
timestamp 1644511149
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_109
timestamp 1644511149
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_121
timestamp 1644511149
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_141
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_153
timestamp 1644511149
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_165
timestamp 1644511149
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_177
timestamp 1644511149
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_189
timestamp 1644511149
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_195
timestamp 1644511149
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_209
timestamp 1644511149
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_221
timestamp 1644511149
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_233
timestamp 1644511149
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_245
timestamp 1644511149
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_251
timestamp 1644511149
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_253
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_267
timestamp 1644511149
transform 1 0 25668 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_279
timestamp 1644511149
transform 1 0 26772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_291
timestamp 1644511149
transform 1 0 27876 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_303
timestamp 1644511149
transform 1 0 28980 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_307
timestamp 1644511149
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_321
timestamp 1644511149
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_333
timestamp 1644511149
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_345
timestamp 1644511149
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_357
timestamp 1644511149
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_363
timestamp 1644511149
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_377
timestamp 1644511149
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_401
timestamp 1644511149
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_413
timestamp 1644511149
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_419
timestamp 1644511149
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_433
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_445
timestamp 1644511149
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_469
timestamp 1644511149
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_475
timestamp 1644511149
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_504
timestamp 1644511149
transform 1 0 47472 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_512
timestamp 1644511149
transform 1 0 48208 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_14
timestamp 1644511149
transform 1 0 2392 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_26
timestamp 1644511149
transform 1 0 3496 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_38
timestamp 1644511149
transform 1 0 4600 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_50
timestamp 1644511149
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_81
timestamp 1644511149
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_93
timestamp 1644511149
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_125
timestamp 1644511149
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_169
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_205
timestamp 1644511149
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_217
timestamp 1644511149
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_223
timestamp 1644511149
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_230
timestamp 1644511149
transform 1 0 22264 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_238
timestamp 1644511149
transform 1 0 23000 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_244
timestamp 1644511149
transform 1 0 23552 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_256
timestamp 1644511149
transform 1 0 24656 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_268
timestamp 1644511149
transform 1 0 25760 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_293
timestamp 1644511149
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_305
timestamp 1644511149
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_317
timestamp 1644511149
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_329
timestamp 1644511149
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_335
timestamp 1644511149
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_373
timestamp 1644511149
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_385
timestamp 1644511149
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_391
timestamp 1644511149
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_393
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_405
timestamp 1644511149
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_417
timestamp 1644511149
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_461
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_473
timestamp 1644511149
transform 1 0 44620 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_485
timestamp 1644511149
transform 1 0 45724 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_497
timestamp 1644511149
transform 1 0 46828 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_505
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_513
timestamp 1644511149
transform 1 0 48300 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_24
timestamp 1644511149
transform 1 0 3312 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_97
timestamp 1644511149
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_109
timestamp 1644511149
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_121
timestamp 1644511149
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_133
timestamp 1644511149
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_141
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_153
timestamp 1644511149
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_177
timestamp 1644511149
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_189
timestamp 1644511149
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_195
timestamp 1644511149
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_200
timestamp 1644511149
transform 1 0 19504 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_204
timestamp 1644511149
transform 1 0 19872 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_213
timestamp 1644511149
transform 1 0 20700 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_239
timestamp 1644511149
transform 1 0 23092 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_248
timestamp 1644511149
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_269
timestamp 1644511149
transform 1 0 25852 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_275
timestamp 1644511149
transform 1 0 26404 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_297
timestamp 1644511149
transform 1 0 28428 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_305
timestamp 1644511149
transform 1 0 29164 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_314
timestamp 1644511149
transform 1 0 29992 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_326
timestamp 1644511149
transform 1 0 31096 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_338
timestamp 1644511149
transform 1 0 32200 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_350
timestamp 1644511149
transform 1 0 33304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_362
timestamp 1644511149
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_377
timestamp 1644511149
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_389
timestamp 1644511149
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_401
timestamp 1644511149
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_413
timestamp 1644511149
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_419
timestamp 1644511149
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_421
timestamp 1644511149
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_433
timestamp 1644511149
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_445
timestamp 1644511149
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_457
timestamp 1644511149
transform 1 0 43148 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_469
timestamp 1644511149
transform 1 0 44252 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_475
timestamp 1644511149
transform 1 0 44804 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_8_489
timestamp 1644511149
transform 1 0 46092 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_8_512
timestamp 1644511149
transform 1 0 48208 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_7
timestamp 1644511149
transform 1 0 1748 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_11
timestamp 1644511149
transform 1 0 2116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_23
timestamp 1644511149
transform 1 0 3220 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_35
timestamp 1644511149
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_47
timestamp 1644511149
transform 1 0 5428 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_57
timestamp 1644511149
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_69
timestamp 1644511149
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_81
timestamp 1644511149
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_93
timestamp 1644511149
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_105
timestamp 1644511149
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_111
timestamp 1644511149
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_113
timestamp 1644511149
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_125
timestamp 1644511149
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_137
timestamp 1644511149
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_149
timestamp 1644511149
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_161
timestamp 1644511149
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_167
timestamp 1644511149
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_169
timestamp 1644511149
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_181
timestamp 1644511149
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_214
timestamp 1644511149
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_222
timestamp 1644511149
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_241
timestamp 1644511149
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_261
timestamp 1644511149
transform 1 0 25116 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_276
timestamp 1644511149
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_309
timestamp 1644511149
transform 1 0 29532 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_331
timestamp 1644511149
transform 1 0 31556 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_335
timestamp 1644511149
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_349
timestamp 1644511149
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_361
timestamp 1644511149
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_385
timestamp 1644511149
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_391
timestamp 1644511149
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_405
timestamp 1644511149
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_429
timestamp 1644511149
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_9_441
timestamp 1644511149
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_447
timestamp 1644511149
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_461
timestamp 1644511149
transform 1 0 43516 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_473
timestamp 1644511149
transform 1 0 44620 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_485
timestamp 1644511149
transform 1 0 45724 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_493
timestamp 1644511149
transform 1 0 46460 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_9_498
timestamp 1644511149
transform 1 0 46920 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_9_508
timestamp 1644511149
transform 1 0 47840 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_13
timestamp 1644511149
transform 1 0 2300 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_25
timestamp 1644511149
transform 1 0 3404 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_10_29
timestamp 1644511149
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_41
timestamp 1644511149
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_53
timestamp 1644511149
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_65
timestamp 1644511149
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_109
timestamp 1644511149
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_141
timestamp 1644511149
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_153
timestamp 1644511149
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_165
timestamp 1644511149
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_177
timestamp 1644511149
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_192
timestamp 1644511149
transform 1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_204
timestamp 1644511149
transform 1 0 19872 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_212
timestamp 1644511149
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_223
timestamp 1644511149
transform 1 0 21620 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_232
timestamp 1644511149
transform 1 0 22448 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_258
timestamp 1644511149
transform 1 0 24840 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_270
timestamp 1644511149
transform 1 0 25944 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_276
timestamp 1644511149
transform 1 0 26496 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_285
timestamp 1644511149
transform 1 0 27324 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_294
timestamp 1644511149
transform 1 0 28152 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_306
timestamp 1644511149
transform 1 0 29256 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_326
timestamp 1644511149
transform 1 0 31096 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_335
timestamp 1644511149
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_347
timestamp 1644511149
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1644511149
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_365
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_377
timestamp 1644511149
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_389
timestamp 1644511149
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_401
timestamp 1644511149
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_413
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_419
timestamp 1644511149
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_421
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_433
timestamp 1644511149
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_445
timestamp 1644511149
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_457
timestamp 1644511149
transform 1 0 43148 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_469
timestamp 1644511149
transform 1 0 44252 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_475
timestamp 1644511149
transform 1 0 44804 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_489
timestamp 1644511149
transform 1 0 46092 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_501
timestamp 1644511149
transform 1 0 47196 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_513
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_3
timestamp 1644511149
transform 1 0 1380 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_25
timestamp 1644511149
transform 1 0 3404 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_37
timestamp 1644511149
transform 1 0 4508 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_49
timestamp 1644511149
transform 1 0 5612 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_57
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_69
timestamp 1644511149
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_81
timestamp 1644511149
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_93
timestamp 1644511149
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_105
timestamp 1644511149
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_111
timestamp 1644511149
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_125
timestamp 1644511149
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_137
timestamp 1644511149
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_149
timestamp 1644511149
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_161
timestamp 1644511149
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_167
timestamp 1644511149
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_11_210
timestamp 1644511149
transform 1 0 20424 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_222
timestamp 1644511149
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_261
timestamp 1644511149
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_273
timestamp 1644511149
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_279
timestamp 1644511149
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_312
timestamp 1644511149
transform 1 0 29808 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_324
timestamp 1644511149
transform 1 0 30912 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_373
timestamp 1644511149
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_385
timestamp 1644511149
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_391
timestamp 1644511149
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_405
timestamp 1644511149
transform 1 0 38364 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_417
timestamp 1644511149
transform 1 0 39468 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_429
timestamp 1644511149
transform 1 0 40572 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_441
timestamp 1644511149
transform 1 0 41676 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_449
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_461
timestamp 1644511149
transform 1 0 43516 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_473
timestamp 1644511149
transform 1 0 44620 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_485
timestamp 1644511149
transform 1 0 45724 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_497
timestamp 1644511149
transform 1 0 46828 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_503
timestamp 1644511149
transform 1 0 47380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_512
timestamp 1644511149
transform 1 0 48208 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_27
timestamp 1644511149
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_29
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_41
timestamp 1644511149
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_53
timestamp 1644511149
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_65
timestamp 1644511149
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_77
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_83
timestamp 1644511149
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_85
timestamp 1644511149
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_97
timestamp 1644511149
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_153
timestamp 1644511149
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_165
timestamp 1644511149
transform 1 0 16284 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_173
timestamp 1644511149
transform 1 0 17020 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_192
timestamp 1644511149
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_208
timestamp 1644511149
transform 1 0 20240 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_228
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_240
timestamp 1644511149
transform 1 0 23184 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_253
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_265
timestamp 1644511149
transform 1 0 25484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_286
timestamp 1644511149
transform 1 0 27416 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_303
timestamp 1644511149
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_307
timestamp 1644511149
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_309
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_321
timestamp 1644511149
transform 1 0 30636 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_333
timestamp 1644511149
transform 1 0 31740 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_357
timestamp 1644511149
transform 1 0 33948 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_365
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_377
timestamp 1644511149
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_389
timestamp 1644511149
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_401
timestamp 1644511149
transform 1 0 37996 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_413
timestamp 1644511149
transform 1 0 39100 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_419
timestamp 1644511149
transform 1 0 39652 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_433
timestamp 1644511149
transform 1 0 40940 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_445
timestamp 1644511149
transform 1 0 42044 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_457
timestamp 1644511149
transform 1 0 43148 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_469
timestamp 1644511149
transform 1 0 44252 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_477
timestamp 1644511149
transform 1 0 44988 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_489
timestamp 1644511149
transform 1 0 46092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_501
timestamp 1644511149
transform 1 0 47196 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_507
timestamp 1644511149
transform 1 0 47748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_512
timestamp 1644511149
transform 1 0 48208 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_27
timestamp 1644511149
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_39
timestamp 1644511149
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_51
timestamp 1644511149
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_55
timestamp 1644511149
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_57
timestamp 1644511149
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_69
timestamp 1644511149
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_81
timestamp 1644511149
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_113
timestamp 1644511149
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_125
timestamp 1644511149
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_137
timestamp 1644511149
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_149
timestamp 1644511149
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_161
timestamp 1644511149
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_167
timestamp 1644511149
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_198
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_215
timestamp 1644511149
transform 1 0 20884 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_223
timestamp 1644511149
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_237
timestamp 1644511149
transform 1 0 22908 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_255
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_276
timestamp 1644511149
transform 1 0 26496 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_289
timestamp 1644511149
transform 1 0 27692 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_13_301
timestamp 1644511149
transform 1 0 28796 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_307
timestamp 1644511149
transform 1 0 29348 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_311
timestamp 1644511149
transform 1 0 29716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_323
timestamp 1644511149
transform 1 0 30820 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_335
timestamp 1644511149
transform 1 0 31924 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_373
timestamp 1644511149
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_385
timestamp 1644511149
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_391
timestamp 1644511149
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_441
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_447
timestamp 1644511149
transform 1 0 42228 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_461
timestamp 1644511149
transform 1 0 43516 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_473
timestamp 1644511149
transform 1 0 44620 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_485
timestamp 1644511149
transform 1 0 45724 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_497
timestamp 1644511149
transform 1 0 46828 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_503
timestamp 1644511149
transform 1 0 47380 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_513
timestamp 1644511149
transform 1 0 48300 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_24
timestamp 1644511149
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_29
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_41
timestamp 1644511149
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_53
timestamp 1644511149
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_65
timestamp 1644511149
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_77
timestamp 1644511149
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_85
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_97
timestamp 1644511149
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_109
timestamp 1644511149
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_121
timestamp 1644511149
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_133
timestamp 1644511149
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_139
timestamp 1644511149
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_141
timestamp 1644511149
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_153
timestamp 1644511149
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_165
timestamp 1644511149
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_177
timestamp 1644511149
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_189
timestamp 1644511149
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_195
timestamp 1644511149
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_202
timestamp 1644511149
transform 1 0 19688 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_216
timestamp 1644511149
transform 1 0 20976 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_228
timestamp 1644511149
transform 1 0 22080 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_236
timestamp 1644511149
transform 1 0 22816 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_248
timestamp 1644511149
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_262
timestamp 1644511149
transform 1 0 25208 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_270
timestamp 1644511149
transform 1 0 25944 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_280
timestamp 1644511149
transform 1 0 26864 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_292
timestamp 1644511149
transform 1 0 27968 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_303
timestamp 1644511149
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_307
timestamp 1644511149
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_314
timestamp 1644511149
transform 1 0 29992 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_336
timestamp 1644511149
transform 1 0 32016 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_348
timestamp 1644511149
transform 1 0 33120 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_360
timestamp 1644511149
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_389
timestamp 1644511149
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_401
timestamp 1644511149
transform 1 0 37996 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_413
timestamp 1644511149
transform 1 0 39100 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_419
timestamp 1644511149
transform 1 0 39652 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_421
timestamp 1644511149
transform 1 0 39836 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_433
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_445
timestamp 1644511149
transform 1 0 42044 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_457
timestamp 1644511149
transform 1 0 43148 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_469
timestamp 1644511149
transform 1 0 44252 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_475
timestamp 1644511149
transform 1 0 44804 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_513
timestamp 1644511149
transform 1 0 48300 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_13
timestamp 1644511149
transform 1 0 2300 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_20
timestamp 1644511149
transform 1 0 2944 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_27
timestamp 1644511149
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_39
timestamp 1644511149
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_51
timestamp 1644511149
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_57
timestamp 1644511149
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_69
timestamp 1644511149
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_81
timestamp 1644511149
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_93
timestamp 1644511149
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_125
timestamp 1644511149
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_137
timestamp 1644511149
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_149
timestamp 1644511149
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_161
timestamp 1644511149
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_193
timestamp 1644511149
transform 1 0 18860 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_15_203
timestamp 1644511149
transform 1 0 19780 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_215
timestamp 1644511149
transform 1 0 20884 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_223
timestamp 1644511149
transform 1 0 21620 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_237
timestamp 1644511149
transform 1 0 22908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_267
timestamp 1644511149
transform 1 0 25668 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_271
timestamp 1644511149
transform 1 0 26036 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_276
timestamp 1644511149
transform 1 0 26496 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_285
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_297
timestamp 1644511149
transform 1 0 28428 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_307
timestamp 1644511149
transform 1 0 29348 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_320
timestamp 1644511149
transform 1 0 30544 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_328
timestamp 1644511149
transform 1 0 31280 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_15_337
timestamp 1644511149
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_349
timestamp 1644511149
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_361
timestamp 1644511149
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_373
timestamp 1644511149
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_385
timestamp 1644511149
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_393
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_405
timestamp 1644511149
transform 1 0 38364 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_417
timestamp 1644511149
transform 1 0 39468 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_429
timestamp 1644511149
transform 1 0 40572 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_441
timestamp 1644511149
transform 1 0 41676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_449
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_461
timestamp 1644511149
transform 1 0 43516 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_473
timestamp 1644511149
transform 1 0 44620 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_485
timestamp 1644511149
transform 1 0 45724 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_500
timestamp 1644511149
transform 1 0 47104 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_512
timestamp 1644511149
transform 1 0 48208 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_24
timestamp 1644511149
transform 1 0 3312 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_29
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_41
timestamp 1644511149
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_53
timestamp 1644511149
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_65
timestamp 1644511149
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_77
timestamp 1644511149
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_83
timestamp 1644511149
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_97
timestamp 1644511149
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_109
timestamp 1644511149
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_121
timestamp 1644511149
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_133
timestamp 1644511149
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_153
timestamp 1644511149
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_165
timestamp 1644511149
transform 1 0 16284 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_16_173
timestamp 1644511149
transform 1 0 17020 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_192
timestamp 1644511149
transform 1 0 18768 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_202
timestamp 1644511149
transform 1 0 19688 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_214
timestamp 1644511149
transform 1 0 20792 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_16_236
timestamp 1644511149
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_248
timestamp 1644511149
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_270
timestamp 1644511149
transform 1 0 25944 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_282
timestamp 1644511149
transform 1 0 27048 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_293
timestamp 1644511149
transform 1 0 28060 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_303
timestamp 1644511149
transform 1 0 28980 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_307
timestamp 1644511149
transform 1 0 29348 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_318
timestamp 1644511149
transform 1 0 30360 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_338
timestamp 1644511149
transform 1 0 32200 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_350
timestamp 1644511149
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_362
timestamp 1644511149
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_365
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_377
timestamp 1644511149
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_389
timestamp 1644511149
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_401
timestamp 1644511149
transform 1 0 37996 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_413
timestamp 1644511149
transform 1 0 39100 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_419
timestamp 1644511149
transform 1 0 39652 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_433
timestamp 1644511149
transform 1 0 40940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_445
timestamp 1644511149
transform 1 0 42044 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_457
timestamp 1644511149
transform 1 0 43148 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_469
timestamp 1644511149
transform 1 0 44252 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_489
timestamp 1644511149
transform 1 0 46092 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_512
timestamp 1644511149
transform 1 0 48208 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_11
timestamp 1644511149
transform 1 0 2116 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_22
timestamp 1644511149
transform 1 0 3128 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_34
timestamp 1644511149
transform 1 0 4232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_17_46
timestamp 1644511149
transform 1 0 5336 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_54
timestamp 1644511149
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_17_57
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_69
timestamp 1644511149
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_93
timestamp 1644511149
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_105
timestamp 1644511149
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_111
timestamp 1644511149
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_125
timestamp 1644511149
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_137
timestamp 1644511149
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_149
timestamp 1644511149
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_161
timestamp 1644511149
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_167
timestamp 1644511149
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_169
timestamp 1644511149
transform 1 0 16652 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_191
timestamp 1644511149
transform 1 0 18676 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_203
timestamp 1644511149
transform 1 0 19780 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_215
timestamp 1644511149
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_223
timestamp 1644511149
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_225
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_229
timestamp 1644511149
transform 1 0 22172 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_241
timestamp 1644511149
transform 1 0 23276 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_247
timestamp 1644511149
transform 1 0 23828 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_257
timestamp 1644511149
transform 1 0 24748 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_265
timestamp 1644511149
transform 1 0 25484 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_276
timestamp 1644511149
transform 1 0 26496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_299
timestamp 1644511149
transform 1 0 28612 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_310
timestamp 1644511149
transform 1 0 29624 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_17_325
timestamp 1644511149
transform 1 0 31004 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_333
timestamp 1644511149
transform 1 0 31740 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_337
timestamp 1644511149
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_349
timestamp 1644511149
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_361
timestamp 1644511149
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_373
timestamp 1644511149
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_385
timestamp 1644511149
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_405
timestamp 1644511149
transform 1 0 38364 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_461
timestamp 1644511149
transform 1 0 43516 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_485
timestamp 1644511149
transform 1 0 45724 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_497
timestamp 1644511149
transform 1 0 46828 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_503
timestamp 1644511149
transform 1 0 47380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_508
timestamp 1644511149
transform 1 0 47840 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_3
timestamp 1644511149
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_15
timestamp 1644511149
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_27
timestamp 1644511149
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_29
timestamp 1644511149
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_41
timestamp 1644511149
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_53
timestamp 1644511149
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_65
timestamp 1644511149
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_77
timestamp 1644511149
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_83
timestamp 1644511149
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_97
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_109
timestamp 1644511149
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_121
timestamp 1644511149
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_133
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_153
timestamp 1644511149
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_165
timestamp 1644511149
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_177
timestamp 1644511149
transform 1 0 17388 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_185
timestamp 1644511149
transform 1 0 18124 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_192
timestamp 1644511149
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_197
timestamp 1644511149
transform 1 0 19228 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_219
timestamp 1644511149
transform 1 0 21252 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_231
timestamp 1644511149
transform 1 0 22356 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_241
timestamp 1644511149
transform 1 0 23276 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_248
timestamp 1644511149
transform 1 0 23920 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_271
timestamp 1644511149
transform 1 0 26036 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_288
timestamp 1644511149
transform 1 0 27600 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_296
timestamp 1644511149
transform 1 0 28336 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_316
timestamp 1644511149
transform 1 0 30176 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_328
timestamp 1644511149
transform 1 0 31280 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_340
timestamp 1644511149
transform 1 0 32384 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_352
timestamp 1644511149
transform 1 0 33488 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_365
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_377
timestamp 1644511149
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_389
timestamp 1644511149
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_401
timestamp 1644511149
transform 1 0 37996 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_413
timestamp 1644511149
transform 1 0 39100 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_419
timestamp 1644511149
transform 1 0 39652 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_433
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_445
timestamp 1644511149
transform 1 0 42044 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_457
timestamp 1644511149
transform 1 0 43148 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_469
timestamp 1644511149
transform 1 0 44252 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_475
timestamp 1644511149
transform 1 0 44804 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_19_13
timestamp 1644511149
transform 1 0 2300 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_25
timestamp 1644511149
transform 1 0 3404 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_37
timestamp 1644511149
transform 1 0 4508 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_49
timestamp 1644511149
transform 1 0 5612 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_55
timestamp 1644511149
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_57
timestamp 1644511149
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_69
timestamp 1644511149
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_81
timestamp 1644511149
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_93
timestamp 1644511149
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_105
timestamp 1644511149
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_111
timestamp 1644511149
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_137
timestamp 1644511149
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_149
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_161
timestamp 1644511149
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_167
timestamp 1644511149
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_169
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_174
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_196
timestamp 1644511149
transform 1 0 19136 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_210
timestamp 1644511149
transform 1 0 20424 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_219
timestamp 1644511149
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_230
timestamp 1644511149
transform 1 0 22264 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_241
timestamp 1644511149
transform 1 0 23276 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_254
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_264
timestamp 1644511149
transform 1 0 25392 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_276
timestamp 1644511149
transform 1 0 26496 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_285
timestamp 1644511149
transform 1 0 27324 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_297
timestamp 1644511149
transform 1 0 28428 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_301
timestamp 1644511149
transform 1 0 28796 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_306
timestamp 1644511149
transform 1 0 29256 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_317
timestamp 1644511149
transform 1 0 30268 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_329
timestamp 1644511149
transform 1 0 31372 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_335
timestamp 1644511149
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_337
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_349
timestamp 1644511149
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_361
timestamp 1644511149
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_373
timestamp 1644511149
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1644511149
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_414
timestamp 1644511149
transform 1 0 39192 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_426
timestamp 1644511149
transform 1 0 40296 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_438
timestamp 1644511149
transform 1 0 41400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_446
timestamp 1644511149
transform 1 0 42136 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_449
timestamp 1644511149
transform 1 0 42412 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_461
timestamp 1644511149
transform 1 0 43516 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_473
timestamp 1644511149
transform 1 0 44620 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_485
timestamp 1644511149
transform 1 0 45724 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_505
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_513
timestamp 1644511149
transform 1 0 48300 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_9
timestamp 1644511149
transform 1 0 1932 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1644511149
transform 1 0 2300 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_25
timestamp 1644511149
transform 1 0 3404 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_53
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_65
timestamp 1644511149
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_77
timestamp 1644511149
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_97
timestamp 1644511149
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_109
timestamp 1644511149
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_121
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_133
timestamp 1644511149
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_139
timestamp 1644511149
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_153
timestamp 1644511149
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_165
timestamp 1644511149
transform 1 0 16284 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_173
timestamp 1644511149
transform 1 0 17020 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_20_178
timestamp 1644511149
transform 1 0 17480 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_190
timestamp 1644511149
transform 1 0 18584 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_213
timestamp 1644511149
transform 1 0 20700 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_225
timestamp 1644511149
transform 1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_245
timestamp 1644511149
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_251
timestamp 1644511149
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_258
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_266
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_274
timestamp 1644511149
transform 1 0 26312 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_286
timestamp 1644511149
transform 1 0 27416 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_294
timestamp 1644511149
transform 1 0 28152 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_20_306
timestamp 1644511149
transform 1 0 29256 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_315
timestamp 1644511149
transform 1 0 30084 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_325
timestamp 1644511149
transform 1 0 31004 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_331
timestamp 1644511149
transform 1 0 31556 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_341
timestamp 1644511149
transform 1 0 32476 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_353
timestamp 1644511149
transform 1 0 33580 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_361
timestamp 1644511149
transform 1 0 34316 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_377
timestamp 1644511149
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_389
timestamp 1644511149
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_401
timestamp 1644511149
transform 1 0 37996 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_413
timestamp 1644511149
transform 1 0 39100 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_419
timestamp 1644511149
transform 1 0 39652 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_433
timestamp 1644511149
transform 1 0 40940 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_445
timestamp 1644511149
transform 1 0 42044 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_457
timestamp 1644511149
transform 1 0 43148 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_469
timestamp 1644511149
transform 1 0 44252 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_475
timestamp 1644511149
transform 1 0 44804 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_477
timestamp 1644511149
transform 1 0 44988 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_489
timestamp 1644511149
transform 1 0 46092 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_501
timestamp 1644511149
transform 1 0 47196 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_513
timestamp 1644511149
transform 1 0 48300 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_28
timestamp 1644511149
transform 1 0 3680 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_40
timestamp 1644511149
transform 1 0 4784 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_52
timestamp 1644511149
transform 1 0 5888 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_81
timestamp 1644511149
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_93
timestamp 1644511149
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_105
timestamp 1644511149
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_113
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_125
timestamp 1644511149
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_137
timestamp 1644511149
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_149
timestamp 1644511149
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_161
timestamp 1644511149
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_167
timestamp 1644511149
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_169
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_173
timestamp 1644511149
transform 1 0 17020 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_195
timestamp 1644511149
transform 1 0 19044 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_206
timestamp 1644511149
transform 1 0 20056 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_215
timestamp 1644511149
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_223
timestamp 1644511149
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_225
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_237
timestamp 1644511149
transform 1 0 22908 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_249
timestamp 1644511149
transform 1 0 24012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_258
timestamp 1644511149
transform 1 0 24840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_266
timestamp 1644511149
transform 1 0 25576 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_276
timestamp 1644511149
transform 1 0 26496 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_285
timestamp 1644511149
transform 1 0 27324 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_294
timestamp 1644511149
transform 1 0 28152 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_21_306
timestamp 1644511149
transform 1 0 29256 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_21_311
timestamp 1644511149
transform 1 0 29716 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_321
timestamp 1644511149
transform 1 0 30636 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_330
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_356
timestamp 1644511149
transform 1 0 33856 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_368
timestamp 1644511149
transform 1 0 34960 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_380
timestamp 1644511149
transform 1 0 36064 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_393
timestamp 1644511149
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_405
timestamp 1644511149
transform 1 0 38364 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_417
timestamp 1644511149
transform 1 0 39468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_429
timestamp 1644511149
transform 1 0 40572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_441
timestamp 1644511149
transform 1 0 41676 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_447
timestamp 1644511149
transform 1 0 42228 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_473
timestamp 1644511149
transform 1 0 44620 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_485
timestamp 1644511149
transform 1 0 45724 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_499
timestamp 1644511149
transform 1 0 47012 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_503
timestamp 1644511149
transform 1 0 47380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_512
timestamp 1644511149
transform 1 0 48208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_3
timestamp 1644511149
transform 1 0 1380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_7
timestamp 1644511149
transform 1 0 1748 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_11
timestamp 1644511149
transform 1 0 2116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_23
timestamp 1644511149
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_27
timestamp 1644511149
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_29
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_41
timestamp 1644511149
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_53
timestamp 1644511149
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_77
timestamp 1644511149
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_97
timestamp 1644511149
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1644511149
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_121
timestamp 1644511149
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_133
timestamp 1644511149
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_139
timestamp 1644511149
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_153
timestamp 1644511149
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_165
timestamp 1644511149
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_177
timestamp 1644511149
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_189
timestamp 1644511149
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_201
timestamp 1644511149
transform 1 0 19596 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_213
timestamp 1644511149
transform 1 0 20700 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_221
timestamp 1644511149
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_239
timestamp 1644511149
transform 1 0 23092 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_251
timestamp 1644511149
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_259
timestamp 1644511149
transform 1 0 24932 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_264
timestamp 1644511149
transform 1 0 25392 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_280
timestamp 1644511149
transform 1 0 26864 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_291
timestamp 1644511149
transform 1 0 27876 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_304
timestamp 1644511149
transform 1 0 29072 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_328
timestamp 1644511149
transform 1 0 31280 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_341
timestamp 1644511149
transform 1 0 32476 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_354
timestamp 1644511149
transform 1 0 33672 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_362
timestamp 1644511149
transform 1 0 34408 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_22_365
timestamp 1644511149
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_377
timestamp 1644511149
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_389
timestamp 1644511149
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_401
timestamp 1644511149
transform 1 0 37996 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_413
timestamp 1644511149
transform 1 0 39100 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_419
timestamp 1644511149
transform 1 0 39652 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_433
timestamp 1644511149
transform 1 0 40940 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_445
timestamp 1644511149
transform 1 0 42044 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_457
timestamp 1644511149
transform 1 0 43148 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_469
timestamp 1644511149
transform 1 0 44252 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_22_489
timestamp 1644511149
transform 1 0 46092 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_512
timestamp 1644511149
transform 1 0 48208 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_15
timestamp 1644511149
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_27
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_39
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_51
timestamp 1644511149
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_55
timestamp 1644511149
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_57
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_69
timestamp 1644511149
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_81
timestamp 1644511149
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_93
timestamp 1644511149
transform 1 0 9660 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_101
timestamp 1644511149
transform 1 0 10396 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_107
timestamp 1644511149
transform 1 0 10948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_111
timestamp 1644511149
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_113
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_125
timestamp 1644511149
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_137
timestamp 1644511149
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_149
timestamp 1644511149
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_161
timestamp 1644511149
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_167
timestamp 1644511149
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_169
timestamp 1644511149
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_181
timestamp 1644511149
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_193
timestamp 1644511149
transform 1 0 18860 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_23_203
timestamp 1644511149
transform 1 0 19780 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_234
timestamp 1644511149
transform 1 0 22632 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_240
timestamp 1644511149
transform 1 0 23184 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_252
timestamp 1644511149
transform 1 0 24288 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_256
timestamp 1644511149
transform 1 0 24656 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_261
timestamp 1644511149
transform 1 0 25116 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_269
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_276
timestamp 1644511149
transform 1 0 26496 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_297
timestamp 1644511149
transform 1 0 28428 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_314
timestamp 1644511149
transform 1 0 29992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_323
timestamp 1644511149
transform 1 0 30820 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_332
timestamp 1644511149
transform 1 0 31648 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_337
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_341
timestamp 1644511149
transform 1 0 32476 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_358
timestamp 1644511149
transform 1 0 34040 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_370
timestamp 1644511149
transform 1 0 35144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_382
timestamp 1644511149
transform 1 0 36248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1644511149
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_405
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_417
timestamp 1644511149
transform 1 0 39468 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_441
timestamp 1644511149
transform 1 0 41676 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_447
timestamp 1644511149
transform 1 0 42228 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_473
timestamp 1644511149
transform 1 0 44620 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_485
timestamp 1644511149
transform 1 0 45724 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_500
timestamp 1644511149
transform 1 0 47104 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_508
timestamp 1644511149
transform 1 0 47840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_29
timestamp 1644511149
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_41
timestamp 1644511149
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_53
timestamp 1644511149
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_65
timestamp 1644511149
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_77
timestamp 1644511149
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_85
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_97
timestamp 1644511149
transform 1 0 10028 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_124
timestamp 1644511149
transform 1 0 12512 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_132
timestamp 1644511149
transform 1 0 13248 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_141
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_153
timestamp 1644511149
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_165
timestamp 1644511149
transform 1 0 16284 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_169
timestamp 1644511149
transform 1 0 16652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1644511149
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_24_197
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_203
timestamp 1644511149
transform 1 0 19780 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_215
timestamp 1644511149
transform 1 0 20884 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_233
timestamp 1644511149
transform 1 0 22540 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_253
timestamp 1644511149
transform 1 0 24380 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_258
timestamp 1644511149
transform 1 0 24840 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_268
timestamp 1644511149
transform 1 0 25760 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_277
timestamp 1644511149
transform 1 0 26588 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_285
timestamp 1644511149
transform 1 0 27324 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_289
timestamp 1644511149
transform 1 0 27692 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_294
timestamp 1644511149
transform 1 0 28152 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_301
timestamp 1644511149
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_307
timestamp 1644511149
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_319
timestamp 1644511149
transform 1 0 30452 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_328
timestamp 1644511149
transform 1 0 31280 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_332
timestamp 1644511149
transform 1 0 31648 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_342
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_354
timestamp 1644511149
transform 1 0 33672 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_362
timestamp 1644511149
transform 1 0 34408 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_421
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_433
timestamp 1644511149
transform 1 0 40940 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_445
timestamp 1644511149
transform 1 0 42044 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_457
timestamp 1644511149
transform 1 0 43148 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_469
timestamp 1644511149
transform 1 0 44252 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_475
timestamp 1644511149
transform 1 0 44804 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_512
timestamp 1644511149
transform 1 0 48208 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_15
timestamp 1644511149
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_27
timestamp 1644511149
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_39
timestamp 1644511149
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_51
timestamp 1644511149
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_55
timestamp 1644511149
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_69
timestamp 1644511149
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_81
timestamp 1644511149
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_93
timestamp 1644511149
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_116
timestamp 1644511149
transform 1 0 11776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_128
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_136
timestamp 1644511149
transform 1 0 13616 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_153
timestamp 1644511149
transform 1 0 15180 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_165
timestamp 1644511149
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_173
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_180
timestamp 1644511149
transform 1 0 17664 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_25_188
timestamp 1644511149
transform 1 0 18400 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_193
timestamp 1644511149
transform 1 0 18860 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_213
timestamp 1644511149
transform 1 0 20700 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_25_221
timestamp 1644511149
transform 1 0 21436 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_228
timestamp 1644511149
transform 1 0 22080 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_239
timestamp 1644511149
transform 1 0 23092 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_250
timestamp 1644511149
transform 1 0 24104 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_254
timestamp 1644511149
transform 1 0 24472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_260
timestamp 1644511149
transform 1 0 25024 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_270
timestamp 1644511149
transform 1 0 25944 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_278
timestamp 1644511149
transform 1 0 26680 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_286
timestamp 1644511149
transform 1 0 27416 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_294
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_298
timestamp 1644511149
transform 1 0 28520 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_304
timestamp 1644511149
transform 1 0 29072 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_315
timestamp 1644511149
transform 1 0 30084 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_328
timestamp 1644511149
transform 1 0 31280 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_343
timestamp 1644511149
transform 1 0 32660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_355
timestamp 1644511149
transform 1 0 33764 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_367
timestamp 1644511149
transform 1 0 34868 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_379
timestamp 1644511149
transform 1 0 35972 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_405
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_417
timestamp 1644511149
transform 1 0 39468 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_429
timestamp 1644511149
transform 1 0 40572 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_441
timestamp 1644511149
transform 1 0 41676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_447
timestamp 1644511149
transform 1 0 42228 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_461
timestamp 1644511149
transform 1 0 43516 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_473
timestamp 1644511149
transform 1 0 44620 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_485
timestamp 1644511149
transform 1 0 45724 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_497
timestamp 1644511149
transform 1 0 46828 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_503
timestamp 1644511149
transform 1 0 47380 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_25_508
timestamp 1644511149
transform 1 0 47840 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_18
timestamp 1644511149
transform 1 0 2760 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_26
timestamp 1644511149
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_32
timestamp 1644511149
transform 1 0 4048 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_44
timestamp 1644511149
transform 1 0 5152 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_56
timestamp 1644511149
transform 1 0 6256 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_80
timestamp 1644511149
transform 1 0 8464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_97
timestamp 1644511149
transform 1 0 10028 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_26_128
timestamp 1644511149
transform 1 0 12880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_151
timestamp 1644511149
transform 1 0 14996 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_172
timestamp 1644511149
transform 1 0 16928 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_179
timestamp 1644511149
transform 1 0 17572 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_187
timestamp 1644511149
transform 1 0 18308 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_192
timestamp 1644511149
transform 1 0 18768 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_202
timestamp 1644511149
transform 1 0 19688 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_210
timestamp 1644511149
transform 1 0 20424 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_26_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_228
timestamp 1644511149
transform 1 0 22080 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_238
timestamp 1644511149
transform 1 0 23000 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_253
timestamp 1644511149
transform 1 0 24380 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_26_265
timestamp 1644511149
transform 1 0 25484 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_279
timestamp 1644511149
transform 1 0 26772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_296
timestamp 1644511149
transform 1 0 28336 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_304
timestamp 1644511149
transform 1 0 29072 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_319
timestamp 1644511149
transform 1 0 30452 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_323
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_340
timestamp 1644511149
transform 1 0 32384 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_353
timestamp 1644511149
transform 1 0 33580 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_361
timestamp 1644511149
transform 1 0 34316 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_26_365
timestamp 1644511149
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_377
timestamp 1644511149
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_389
timestamp 1644511149
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_401
timestamp 1644511149
transform 1 0 37996 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_457
timestamp 1644511149
transform 1 0 43148 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_469
timestamp 1644511149
transform 1 0 44252 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_489
timestamp 1644511149
transform 1 0 46092 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_512
timestamp 1644511149
transform 1 0 48208 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_24
timestamp 1644511149
transform 1 0 3312 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_69
timestamp 1644511149
transform 1 0 7452 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_89
timestamp 1644511149
transform 1 0 9292 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_101
timestamp 1644511149
transform 1 0 10396 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_109
timestamp 1644511149
transform 1 0 11132 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_27_147
timestamp 1644511149
transform 1 0 14628 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_173
timestamp 1644511149
transform 1 0 17020 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_180
timestamp 1644511149
transform 1 0 17664 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_200
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_27_210
timestamp 1644511149
transform 1 0 20424 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_222
timestamp 1644511149
transform 1 0 21528 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_229
timestamp 1644511149
transform 1 0 22172 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_241
timestamp 1644511149
transform 1 0 23276 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_250
timestamp 1644511149
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_27_254
timestamp 1644511149
transform 1 0 24472 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_27_262
timestamp 1644511149
transform 1 0 25208 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_270
timestamp 1644511149
transform 1 0 25944 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_276
timestamp 1644511149
transform 1 0 26496 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_285
timestamp 1644511149
transform 1 0 27324 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_296
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_306
timestamp 1644511149
transform 1 0 29256 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_319
timestamp 1644511149
transform 1 0 30452 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_331
timestamp 1644511149
transform 1 0 31556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_335
timestamp 1644511149
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_353
timestamp 1644511149
transform 1 0 33580 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_365
timestamp 1644511149
transform 1 0 34684 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_377
timestamp 1644511149
transform 1 0 35788 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_389
timestamp 1644511149
transform 1 0 36892 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_27_393
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_405
timestamp 1644511149
transform 1 0 38364 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_417
timestamp 1644511149
transform 1 0 39468 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_429
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_441
timestamp 1644511149
transform 1 0 41676 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_447
timestamp 1644511149
transform 1 0 42228 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_500
timestamp 1644511149
transform 1 0 47104 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_508
timestamp 1644511149
transform 1 0 47840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_24
timestamp 1644511149
transform 1 0 3312 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_53
timestamp 1644511149
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_65
timestamp 1644511149
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_71
timestamp 1644511149
transform 1 0 7636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_80
timestamp 1644511149
transform 1 0 8464 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_93
timestamp 1644511149
transform 1 0 9660 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_101
timestamp 1644511149
transform 1 0 10396 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_120
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_128
timestamp 1644511149
transform 1 0 12880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_136
timestamp 1644511149
transform 1 0 13616 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_161
timestamp 1644511149
transform 1 0 15916 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_169
timestamp 1644511149
transform 1 0 16652 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_175
timestamp 1644511149
transform 1 0 17204 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_180
timestamp 1644511149
transform 1 0 17664 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_192
timestamp 1644511149
transform 1 0 18768 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_213
timestamp 1644511149
transform 1 0 20700 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_221
timestamp 1644511149
transform 1 0 21436 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_242
timestamp 1644511149
transform 1 0 23368 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_250
timestamp 1644511149
transform 1 0 24104 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_28_253
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_266
timestamp 1644511149
transform 1 0 25576 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_273
timestamp 1644511149
transform 1 0 26220 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_281
timestamp 1644511149
transform 1 0 26956 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_293
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_301
timestamp 1644511149
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_315
timestamp 1644511149
transform 1 0 30084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_327
timestamp 1644511149
transform 1 0 31188 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_339
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_351
timestamp 1644511149
transform 1 0 33396 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_363
timestamp 1644511149
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_389
timestamp 1644511149
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_401
timestamp 1644511149
transform 1 0 37996 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_413
timestamp 1644511149
transform 1 0 39100 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_419
timestamp 1644511149
transform 1 0 39652 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_433
timestamp 1644511149
transform 1 0 40940 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_445
timestamp 1644511149
transform 1 0 42044 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_457
timestamp 1644511149
transform 1 0 43148 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_469
timestamp 1644511149
transform 1 0 44252 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_475
timestamp 1644511149
transform 1 0 44804 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_477
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_489
timestamp 1644511149
transform 1 0 46092 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_28_501
timestamp 1644511149
transform 1 0 47196 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_515
timestamp 1644511149
transform 1 0 48484 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_6
timestamp 1644511149
transform 1 0 1656 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_20
timestamp 1644511149
transform 1 0 2944 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_32
timestamp 1644511149
transform 1 0 4048 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_44
timestamp 1644511149
transform 1 0 5152 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_69
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_89
timestamp 1644511149
transform 1 0 9292 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_101
timestamp 1644511149
transform 1 0 10396 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_29_113
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_124
timestamp 1644511149
transform 1 0 12512 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_132
timestamp 1644511149
transform 1 0 13248 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_142
timestamp 1644511149
transform 1 0 14168 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_150
timestamp 1644511149
transform 1 0 14904 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_154
timestamp 1644511149
transform 1 0 15272 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_159
timestamp 1644511149
transform 1 0 15732 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_167
timestamp 1644511149
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_173
timestamp 1644511149
transform 1 0 17020 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_181
timestamp 1644511149
transform 1 0 17756 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_191
timestamp 1644511149
transform 1 0 18676 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_195
timestamp 1644511149
transform 1 0 19044 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_201
timestamp 1644511149
transform 1 0 19596 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_213
timestamp 1644511149
transform 1 0 20700 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_221
timestamp 1644511149
transform 1 0 21436 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_241
timestamp 1644511149
transform 1 0 23276 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_250
timestamp 1644511149
transform 1 0 24104 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_256
timestamp 1644511149
transform 1 0 24656 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_262
timestamp 1644511149
transform 1 0 25208 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_275
timestamp 1644511149
transform 1 0 26404 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_279
timestamp 1644511149
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_281
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_287
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_304
timestamp 1644511149
transform 1 0 29072 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_316
timestamp 1644511149
transform 1 0 30176 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_328
timestamp 1644511149
transform 1 0 31280 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_29_337
timestamp 1644511149
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_349
timestamp 1644511149
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_361
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_373
timestamp 1644511149
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_385
timestamp 1644511149
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_391
timestamp 1644511149
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_393
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_405
timestamp 1644511149
transform 1 0 38364 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_429
timestamp 1644511149
transform 1 0 40572 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_441
timestamp 1644511149
transform 1 0 41676 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_473
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_485
timestamp 1644511149
transform 1 0 45724 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_497
timestamp 1644511149
transform 1 0 46828 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_503
timestamp 1644511149
transform 1 0 47380 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_513
timestamp 1644511149
transform 1 0 48300 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1644511149
transform 1 0 1380 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_15
timestamp 1644511149
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_27
timestamp 1644511149
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_29
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_41
timestamp 1644511149
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_53
timestamp 1644511149
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_68
timestamp 1644511149
transform 1 0 7360 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_74
timestamp 1644511149
transform 1 0 7912 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_78
timestamp 1644511149
transform 1 0 8280 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_30_93
timestamp 1644511149
transform 1 0 9660 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_117
timestamp 1644511149
transform 1 0 11868 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_131
timestamp 1644511149
transform 1 0 13156 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_139
timestamp 1644511149
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_153
timestamp 1644511149
transform 1 0 15180 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_30_169
timestamp 1644511149
transform 1 0 16652 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_192
timestamp 1644511149
transform 1 0 18768 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_197
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_209
timestamp 1644511149
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_221
timestamp 1644511149
transform 1 0 21436 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_229
timestamp 1644511149
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_236
timestamp 1644511149
transform 1 0 22816 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_253
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_266
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_277
timestamp 1644511149
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_30_295
timestamp 1644511149
transform 1 0 28244 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_309
timestamp 1644511149
transform 1 0 29532 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_317
timestamp 1644511149
transform 1 0 30268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_329
timestamp 1644511149
transform 1 0 31372 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_339
timestamp 1644511149
transform 1 0 32292 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_351
timestamp 1644511149
transform 1 0 33396 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_363
timestamp 1644511149
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_389
timestamp 1644511149
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_401
timestamp 1644511149
transform 1 0 37996 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_413
timestamp 1644511149
transform 1 0 39100 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_433
timestamp 1644511149
transform 1 0 40940 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_445
timestamp 1644511149
transform 1 0 42044 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_457
timestamp 1644511149
transform 1 0 43148 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_469
timestamp 1644511149
transform 1 0 44252 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_475
timestamp 1644511149
transform 1 0 44804 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_512
timestamp 1644511149
transform 1 0 48208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_3
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_7
timestamp 1644511149
transform 1 0 1748 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_29
timestamp 1644511149
transform 1 0 3772 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_41
timestamp 1644511149
transform 1 0 4876 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_53
timestamp 1644511149
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_69
timestamp 1644511149
transform 1 0 7452 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_93
timestamp 1644511149
transform 1 0 9660 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_101
timestamp 1644511149
transform 1 0 10396 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_108
timestamp 1644511149
transform 1 0 11040 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_31_127
timestamp 1644511149
transform 1 0 12788 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_147
timestamp 1644511149
transform 1 0 14628 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_159
timestamp 1644511149
transform 1 0 15732 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1644511149
transform 1 0 16192 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_169
timestamp 1644511149
transform 1 0 16652 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_186
timestamp 1644511149
transform 1 0 18216 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_194
timestamp 1644511149
transform 1 0 18952 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_202
timestamp 1644511149
transform 1 0 19688 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_208
timestamp 1644511149
transform 1 0 20240 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_225
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_233
timestamp 1644511149
transform 1 0 22540 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_237
timestamp 1644511149
transform 1 0 22908 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_259
timestamp 1644511149
transform 1 0 24932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_267
timestamp 1644511149
transform 1 0 25668 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_274
timestamp 1644511149
transform 1 0 26312 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_293
timestamp 1644511149
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_307
timestamp 1644511149
transform 1 0 29348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_315
timestamp 1644511149
transform 1 0 30084 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_31_325
timestamp 1644511149
transform 1 0 31004 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_333
timestamp 1644511149
transform 1 0 31740 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_31_337
timestamp 1644511149
transform 1 0 32108 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_354
timestamp 1644511149
transform 1 0 33672 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_366
timestamp 1644511149
transform 1 0 34776 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_378
timestamp 1644511149
transform 1 0 35880 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_390
timestamp 1644511149
transform 1 0 36984 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_405
timestamp 1644511149
transform 1 0 38364 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_417
timestamp 1644511149
transform 1 0 39468 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_429
timestamp 1644511149
transform 1 0 40572 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_31_441
timestamp 1644511149
transform 1 0 41676 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_447
timestamp 1644511149
transform 1 0 42228 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_461
timestamp 1644511149
transform 1 0 43516 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_473
timestamp 1644511149
transform 1 0 44620 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_485
timestamp 1644511149
transform 1 0 45724 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_493
timestamp 1644511149
transform 1 0 46460 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_31_498
timestamp 1644511149
transform 1 0 46920 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_508
timestamp 1644511149
transform 1 0 47840 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_7
timestamp 1644511149
transform 1 0 1748 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_11
timestamp 1644511149
transform 1 0 2116 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_23
timestamp 1644511149
transform 1 0 3220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_27
timestamp 1644511149
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_41
timestamp 1644511149
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_53
timestamp 1644511149
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_65
timestamp 1644511149
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_77
timestamp 1644511149
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_83
timestamp 1644511149
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_97
timestamp 1644511149
transform 1 0 10028 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_114
timestamp 1644511149
transform 1 0 11592 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_123
timestamp 1644511149
transform 1 0 12420 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_146
timestamp 1644511149
transform 1 0 14536 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_158
timestamp 1644511149
transform 1 0 15640 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_166
timestamp 1644511149
transform 1 0 16376 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_32_177
timestamp 1644511149
transform 1 0 17388 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_183
timestamp 1644511149
transform 1 0 17940 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_192
timestamp 1644511149
transform 1 0 18768 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_214
timestamp 1644511149
transform 1 0 20792 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_234
timestamp 1644511149
transform 1 0 22632 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_246
timestamp 1644511149
transform 1 0 23736 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_269
timestamp 1644511149
transform 1 0 25852 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_277
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_293
timestamp 1644511149
transform 1 0 28060 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_305
timestamp 1644511149
transform 1 0 29164 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_325
timestamp 1644511149
transform 1 0 31004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_334
timestamp 1644511149
transform 1 0 31832 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_343
timestamp 1644511149
transform 1 0 32660 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_351
timestamp 1644511149
transform 1 0 33396 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_359
timestamp 1644511149
transform 1 0 34132 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_363
timestamp 1644511149
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_381
timestamp 1644511149
transform 1 0 36156 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_393
timestamp 1644511149
transform 1 0 37260 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_405
timestamp 1644511149
transform 1 0 38364 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_417
timestamp 1644511149
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_457
timestamp 1644511149
transform 1 0 43148 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_32_469
timestamp 1644511149
transform 1 0 44252 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_475
timestamp 1644511149
transform 1 0 44804 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_32_512
timestamp 1644511149
transform 1 0 48208 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1644511149
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_27
timestamp 1644511149
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_39
timestamp 1644511149
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_51
timestamp 1644511149
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_55
timestamp 1644511149
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_60
timestamp 1644511149
transform 1 0 6624 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_84
timestamp 1644511149
transform 1 0 8832 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_93
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_101
timestamp 1644511149
transform 1 0 10396 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_108
timestamp 1644511149
transform 1 0 11040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_117
timestamp 1644511149
transform 1 0 11868 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_33_126
timestamp 1644511149
transform 1 0 12696 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_132
timestamp 1644511149
transform 1 0 13248 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_141
timestamp 1644511149
transform 1 0 14076 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1644511149
transform 1 0 15180 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_163
timestamp 1644511149
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_167
timestamp 1644511149
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_177
timestamp 1644511149
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_189
timestamp 1644511149
transform 1 0 18492 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_197
timestamp 1644511149
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_204
timestamp 1644511149
transform 1 0 19872 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_216
timestamp 1644511149
transform 1 0 20976 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_225
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_237
timestamp 1644511149
transform 1 0 22908 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_244
timestamp 1644511149
transform 1 0 23552 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_256
timestamp 1644511149
transform 1 0 24656 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_268
timestamp 1644511149
transform 1 0 25760 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_281
timestamp 1644511149
transform 1 0 26956 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_289
timestamp 1644511149
transform 1 0 27692 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_295
timestamp 1644511149
transform 1 0 28244 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_307
timestamp 1644511149
transform 1 0 29348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_315
timestamp 1644511149
transform 1 0 30084 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_332
timestamp 1644511149
transform 1 0 31648 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_353
timestamp 1644511149
transform 1 0 33580 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_365
timestamp 1644511149
transform 1 0 34684 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_377
timestamp 1644511149
transform 1 0 35788 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1644511149
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_405
timestamp 1644511149
transform 1 0 38364 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_417
timestamp 1644511149
transform 1 0 39468 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_429
timestamp 1644511149
transform 1 0 40572 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_441
timestamp 1644511149
transform 1 0 41676 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_447
timestamp 1644511149
transform 1 0 42228 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_449
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_461
timestamp 1644511149
transform 1 0 43516 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_473
timestamp 1644511149
transform 1 0 44620 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_485
timestamp 1644511149
transform 1 0 45724 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_497
timestamp 1644511149
transform 1 0 46828 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_503
timestamp 1644511149
transform 1 0 47380 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_513
timestamp 1644511149
transform 1 0 48300 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1644511149
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_27
timestamp 1644511149
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_34_77
timestamp 1644511149
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_83
timestamp 1644511149
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_93
timestamp 1644511149
transform 1 0 9660 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_34_122
timestamp 1644511149
transform 1 0 12328 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_134
timestamp 1644511149
transform 1 0 13432 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_34_141
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_159
timestamp 1644511149
transform 1 0 15732 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_179
timestamp 1644511149
transform 1 0 17572 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_191
timestamp 1644511149
transform 1 0 18676 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_195
timestamp 1644511149
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_197
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_205
timestamp 1644511149
transform 1 0 19964 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_211
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_216
timestamp 1644511149
transform 1 0 20976 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_228
timestamp 1644511149
transform 1 0 22080 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_236
timestamp 1644511149
transform 1 0 22816 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_258
timestamp 1644511149
transform 1 0 24840 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_270
timestamp 1644511149
transform 1 0 25944 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_276
timestamp 1644511149
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_307
timestamp 1644511149
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_309
timestamp 1644511149
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_321
timestamp 1644511149
transform 1 0 30636 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_327
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_336
timestamp 1644511149
transform 1 0 32016 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_345
timestamp 1644511149
transform 1 0 32844 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_34_358
timestamp 1644511149
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_34_365
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_377
timestamp 1644511149
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_389
timestamp 1644511149
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_401
timestamp 1644511149
transform 1 0 37996 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_413
timestamp 1644511149
transform 1 0 39100 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_433
timestamp 1644511149
transform 1 0 40940 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_445
timestamp 1644511149
transform 1 0 42044 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_457
timestamp 1644511149
transform 1 0 43148 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_469
timestamp 1644511149
transform 1 0 44252 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_477
timestamp 1644511149
transform 1 0 44988 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_489
timestamp 1644511149
transform 1 0 46092 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_501
timestamp 1644511149
transform 1 0 47196 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_513
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_3
timestamp 1644511149
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_15
timestamp 1644511149
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_27
timestamp 1644511149
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_39
timestamp 1644511149
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_51
timestamp 1644511149
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_55
timestamp 1644511149
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_85
timestamp 1644511149
transform 1 0 8924 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_97
timestamp 1644511149
transform 1 0 10028 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_109
timestamp 1644511149
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_116
timestamp 1644511149
transform 1 0 11776 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_35_128
timestamp 1644511149
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1644511149
transform 1 0 13616 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_150
timestamp 1644511149
transform 1 0 14904 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_162
timestamp 1644511149
transform 1 0 16008 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_185
timestamp 1644511149
transform 1 0 18124 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_193
timestamp 1644511149
transform 1 0 18860 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_199
timestamp 1644511149
transform 1 0 19412 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_206
timestamp 1644511149
transform 1 0 20056 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_216
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_244
timestamp 1644511149
transform 1 0 23552 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_258
timestamp 1644511149
transform 1 0 24840 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_35_272
timestamp 1644511149
transform 1 0 26128 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_35_286
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_294
timestamp 1644511149
transform 1 0 28152 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_303
timestamp 1644511149
transform 1 0 28980 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_312
timestamp 1644511149
transform 1 0 29808 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_321
timestamp 1644511149
transform 1 0 30636 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_333
timestamp 1644511149
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_349
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_371
timestamp 1644511149
transform 1 0 35236 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_35_383
timestamp 1644511149
transform 1 0 36340 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_391
timestamp 1644511149
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_461
timestamp 1644511149
transform 1 0 43516 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_473
timestamp 1644511149
transform 1 0 44620 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_485
timestamp 1644511149
transform 1 0 45724 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_497
timestamp 1644511149
transform 1 0 46828 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_35_512
timestamp 1644511149
transform 1 0 48208 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_15
timestamp 1644511149
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_27
timestamp 1644511149
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_41
timestamp 1644511149
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_53
timestamp 1644511149
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_65
timestamp 1644511149
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_77
timestamp 1644511149
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_83
timestamp 1644511149
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_36_90
timestamp 1644511149
transform 1 0 9384 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_98
timestamp 1644511149
transform 1 0 10120 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_102
timestamp 1644511149
transform 1 0 10488 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_127
timestamp 1644511149
transform 1 0 12788 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_139
timestamp 1644511149
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_146
timestamp 1644511149
transform 1 0 14536 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_158
timestamp 1644511149
transform 1 0 15640 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_170
timestamp 1644511149
transform 1 0 16744 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_182
timestamp 1644511149
transform 1 0 17848 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_192
timestamp 1644511149
transform 1 0 18768 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_213
timestamp 1644511149
transform 1 0 20700 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_217
timestamp 1644511149
transform 1 0 21068 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_226
timestamp 1644511149
transform 1 0 21896 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_238
timestamp 1644511149
transform 1 0 23000 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_244
timestamp 1644511149
transform 1 0 23552 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_259
timestamp 1644511149
transform 1 0 24932 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_265
timestamp 1644511149
transform 1 0 25484 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_36_282
timestamp 1644511149
transform 1 0 27048 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_330
timestamp 1644511149
transform 1 0 31464 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_342
timestamp 1644511149
transform 1 0 32568 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_348
timestamp 1644511149
transform 1 0 33120 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_381
timestamp 1644511149
transform 1 0 36156 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_393
timestamp 1644511149
transform 1 0 37260 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_405
timestamp 1644511149
transform 1 0 38364 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_417
timestamp 1644511149
transform 1 0 39468 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_433
timestamp 1644511149
transform 1 0 40940 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_445
timestamp 1644511149
transform 1 0 42044 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_457
timestamp 1644511149
transform 1 0 43148 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_469
timestamp 1644511149
transform 1 0 44252 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_475
timestamp 1644511149
transform 1 0 44804 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_489
timestamp 1644511149
transform 1 0 46092 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_36_501
timestamp 1644511149
transform 1 0 47196 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_512
timestamp 1644511149
transform 1 0 48208 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_11
timestamp 1644511149
transform 1 0 2116 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_18
timestamp 1644511149
transform 1 0 2760 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_30
timestamp 1644511149
transform 1 0 3864 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_42
timestamp 1644511149
transform 1 0 4968 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_37_54
timestamp 1644511149
transform 1 0 6072 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_81
timestamp 1644511149
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_93
timestamp 1644511149
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_105
timestamp 1644511149
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_111
timestamp 1644511149
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_113
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_125
timestamp 1644511149
transform 1 0 12604 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_129
timestamp 1644511149
transform 1 0 12972 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_137
timestamp 1644511149
transform 1 0 13708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_145
timestamp 1644511149
transform 1 0 14444 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_157
timestamp 1644511149
transform 1 0 15548 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_165
timestamp 1644511149
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_173
timestamp 1644511149
transform 1 0 17020 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_193
timestamp 1644511149
transform 1 0 18860 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_207
timestamp 1644511149
transform 1 0 20148 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_216
timestamp 1644511149
transform 1 0 20976 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_242
timestamp 1644511149
transform 1 0 23368 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_249
timestamp 1644511149
transform 1 0 24012 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_257
timestamp 1644511149
transform 1 0 24748 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_37_264
timestamp 1644511149
transform 1 0 25392 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_270
timestamp 1644511149
transform 1 0 25944 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_291
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_303
timestamp 1644511149
transform 1 0 28980 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_312
timestamp 1644511149
transform 1 0 29808 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_332
timestamp 1644511149
transform 1 0 31648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_349
timestamp 1644511149
transform 1 0 33212 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_363
timestamp 1644511149
transform 1 0 34500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_375
timestamp 1644511149
transform 1 0 35604 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_387
timestamp 1644511149
transform 1 0 36708 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_391
timestamp 1644511149
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_393
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_405
timestamp 1644511149
transform 1 0 38364 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_417
timestamp 1644511149
transform 1 0 39468 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_429
timestamp 1644511149
transform 1 0 40572 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_441
timestamp 1644511149
transform 1 0 41676 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_447
timestamp 1644511149
transform 1 0 42228 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_461
timestamp 1644511149
transform 1 0 43516 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_473
timestamp 1644511149
transform 1 0 44620 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_485
timestamp 1644511149
transform 1 0 45724 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_497
timestamp 1644511149
transform 1 0 46828 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_503
timestamp 1644511149
transform 1 0 47380 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_512
timestamp 1644511149
transform 1 0 48208 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_24
timestamp 1644511149
transform 1 0 3312 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_41
timestamp 1644511149
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_53
timestamp 1644511149
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_65
timestamp 1644511149
transform 1 0 7084 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_71
timestamp 1644511149
transform 1 0 7636 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_75
timestamp 1644511149
transform 1 0 8004 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_83
timestamp 1644511149
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_94
timestamp 1644511149
transform 1 0 9752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_117
timestamp 1644511149
transform 1 0 11868 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_123
timestamp 1644511149
transform 1 0 12420 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_130
timestamp 1644511149
transform 1 0 13064 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_138
timestamp 1644511149
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_38_146
timestamp 1644511149
transform 1 0 14536 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_154
timestamp 1644511149
transform 1 0 15272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_38_174
timestamp 1644511149
transform 1 0 17112 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_185
timestamp 1644511149
transform 1 0 18124 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_193
timestamp 1644511149
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_205
timestamp 1644511149
transform 1 0 19964 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_220
timestamp 1644511149
transform 1 0 21344 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_232
timestamp 1644511149
transform 1 0 22448 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_244
timestamp 1644511149
transform 1 0 23552 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_259
timestamp 1644511149
transform 1 0 24932 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_267
timestamp 1644511149
transform 1 0 25668 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_279
timestamp 1644511149
transform 1 0 26772 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_291
timestamp 1644511149
transform 1 0 27876 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_38_302
timestamp 1644511149
transform 1 0 28888 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_38_309
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_321
timestamp 1644511149
transform 1 0 30636 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_328
timestamp 1644511149
transform 1 0 31280 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_340
timestamp 1644511149
transform 1 0 32384 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_352
timestamp 1644511149
transform 1 0 33488 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_489
timestamp 1644511149
transform 1 0 46092 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_501
timestamp 1644511149
transform 1 0 47196 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_38_513
timestamp 1644511149
transform 1 0 48300 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_7
timestamp 1644511149
transform 1 0 1748 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_11
timestamp 1644511149
transform 1 0 2116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_23
timestamp 1644511149
transform 1 0 3220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_35
timestamp 1644511149
transform 1 0 4324 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_47
timestamp 1644511149
transform 1 0 5428 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_55
timestamp 1644511149
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_65
timestamp 1644511149
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_89
timestamp 1644511149
transform 1 0 9292 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_97
timestamp 1644511149
transform 1 0 10028 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_109
timestamp 1644511149
transform 1 0 11132 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_120
timestamp 1644511149
transform 1 0 12144 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_128
timestamp 1644511149
transform 1 0 12880 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1644511149
transform 1 0 13892 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_149
timestamp 1644511149
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_161
timestamp 1644511149
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_167
timestamp 1644511149
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_177
timestamp 1644511149
transform 1 0 17388 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_181
timestamp 1644511149
transform 1 0 17756 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_190
timestamp 1644511149
transform 1 0 18584 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_196
timestamp 1644511149
transform 1 0 19136 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_202
timestamp 1644511149
transform 1 0 19688 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_208
timestamp 1644511149
transform 1 0 20240 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_244
timestamp 1644511149
transform 1 0 23552 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_258
timestamp 1644511149
transform 1 0 24840 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_266
timestamp 1644511149
transform 1 0 25576 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_276
timestamp 1644511149
transform 1 0 26496 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_286
timestamp 1644511149
transform 1 0 27416 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_290
timestamp 1644511149
transform 1 0 27784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_299
timestamp 1644511149
transform 1 0 28612 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_332
timestamp 1644511149
transform 1 0 31648 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_341
timestamp 1644511149
transform 1 0 32476 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_345
timestamp 1644511149
transform 1 0 32844 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_370
timestamp 1644511149
transform 1 0 35144 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_382
timestamp 1644511149
transform 1 0 36248 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_390
timestamp 1644511149
transform 1 0 36984 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_393
timestamp 1644511149
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_405
timestamp 1644511149
transform 1 0 38364 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_417
timestamp 1644511149
transform 1 0 39468 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_473
timestamp 1644511149
transform 1 0 44620 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_485
timestamp 1644511149
transform 1 0 45724 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_497
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_503
timestamp 1644511149
transform 1 0 47380 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_39_505
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_512
timestamp 1644511149
transform 1 0 48208 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_7
timestamp 1644511149
transform 1 0 1748 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_19
timestamp 1644511149
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_29
timestamp 1644511149
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_41
timestamp 1644511149
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_53
timestamp 1644511149
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_65
timestamp 1644511149
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_40_77
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_103
timestamp 1644511149
transform 1 0 10580 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_115
timestamp 1644511149
transform 1 0 11684 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_123
timestamp 1644511149
transform 1 0 12420 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_40_131
timestamp 1644511149
transform 1 0 13156 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_139
timestamp 1644511149
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_141
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_153
timestamp 1644511149
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_165
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_171
timestamp 1644511149
transform 1 0 16836 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_183
timestamp 1644511149
transform 1 0 17940 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_201
timestamp 1644511149
transform 1 0 19596 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_219
timestamp 1644511149
transform 1 0 21252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_243
timestamp 1644511149
transform 1 0 23460 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_251
timestamp 1644511149
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_40_259
timestamp 1644511149
transform 1 0 24932 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_267
timestamp 1644511149
transform 1 0 25668 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_284
timestamp 1644511149
transform 1 0 27232 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_304
timestamp 1644511149
transform 1 0 29072 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_318
timestamp 1644511149
transform 1 0 30360 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_325
timestamp 1644511149
transform 1 0 31004 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_350
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_357
timestamp 1644511149
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_386
timestamp 1644511149
transform 1 0 36616 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_398
timestamp 1644511149
transform 1 0 37720 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_410
timestamp 1644511149
transform 1 0 38824 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_418
timestamp 1644511149
transform 1 0 39560 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_427
timestamp 1644511149
transform 1 0 40388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_439
timestamp 1644511149
transform 1 0 41492 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_451
timestamp 1644511149
transform 1 0 42596 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_463
timestamp 1644511149
transform 1 0 43700 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_475
timestamp 1644511149
transform 1 0 44804 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_477
timestamp 1644511149
transform 1 0 44988 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_489
timestamp 1644511149
transform 1 0 46092 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_512
timestamp 1644511149
transform 1 0 48208 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_15
timestamp 1644511149
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_27
timestamp 1644511149
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_39
timestamp 1644511149
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_51
timestamp 1644511149
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_55
timestamp 1644511149
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_69
timestamp 1644511149
transform 1 0 7452 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_75
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_85
timestamp 1644511149
transform 1 0 8924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_97
timestamp 1644511149
transform 1 0 10028 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_108
timestamp 1644511149
transform 1 0 11040 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_133
timestamp 1644511149
transform 1 0 13340 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_138
timestamp 1644511149
transform 1 0 13800 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_150
timestamp 1644511149
transform 1 0 14904 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_162
timestamp 1644511149
transform 1 0 16008 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_181
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_193
timestamp 1644511149
transform 1 0 18860 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_199
timestamp 1644511149
transform 1 0 19412 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_41_207
timestamp 1644511149
transform 1 0 20148 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_41_218
timestamp 1644511149
transform 1 0 21160 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_233
timestamp 1644511149
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_41_236
timestamp 1644511149
transform 1 0 22816 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_244
timestamp 1644511149
transform 1 0 23552 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_254
timestamp 1644511149
transform 1 0 24472 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_262
timestamp 1644511149
transform 1 0 25208 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_266
timestamp 1644511149
transform 1 0 25576 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_274
timestamp 1644511149
transform 1 0 26312 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_41_285
timestamp 1644511149
transform 1 0 27324 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_291
timestamp 1644511149
transform 1 0 27876 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_298
timestamp 1644511149
transform 1 0 28520 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_41_314
timestamp 1644511149
transform 1 0 29992 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_332
timestamp 1644511149
transform 1 0 31648 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_340
timestamp 1644511149
transform 1 0 32384 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_365
timestamp 1644511149
transform 1 0 34684 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_377
timestamp 1644511149
transform 1 0 35788 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_389
timestamp 1644511149
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_408
timestamp 1644511149
transform 1 0 38640 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_420
timestamp 1644511149
transform 1 0 39744 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_41_444
timestamp 1644511149
transform 1 0 41952 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_473
timestamp 1644511149
transform 1 0 44620 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_485
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_500
timestamp 1644511149
transform 1 0 47104 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_508
timestamp 1644511149
transform 1 0 47840 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_15
timestamp 1644511149
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_27
timestamp 1644511149
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_29
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_41
timestamp 1644511149
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_53
timestamp 1644511149
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_65
timestamp 1644511149
transform 1 0 7084 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_73
timestamp 1644511149
transform 1 0 7820 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_80
timestamp 1644511149
transform 1 0 8464 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_96
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_107
timestamp 1644511149
transform 1 0 10948 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_115
timestamp 1644511149
transform 1 0 11684 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_123
timestamp 1644511149
transform 1 0 12420 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_147
timestamp 1644511149
transform 1 0 14628 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_159
timestamp 1644511149
transform 1 0 15732 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_163
timestamp 1644511149
transform 1 0 16100 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_180
timestamp 1644511149
transform 1 0 17664 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_192
timestamp 1644511149
transform 1 0 18768 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_207
timestamp 1644511149
transform 1 0 20148 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_227
timestamp 1644511149
transform 1 0 21988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_245
timestamp 1644511149
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_42_253
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_259
timestamp 1644511149
transform 1 0 24932 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_267
timestamp 1644511149
transform 1 0 25668 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_287
timestamp 1644511149
transform 1 0 27508 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_333
timestamp 1644511149
transform 1 0 31740 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_349
timestamp 1644511149
transform 1 0 33212 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_357
timestamp 1644511149
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_363
timestamp 1644511149
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_368
timestamp 1644511149
transform 1 0 34960 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_380
timestamp 1644511149
transform 1 0 36064 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_392
timestamp 1644511149
transform 1 0 37168 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_404
timestamp 1644511149
transform 1 0 38272 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_416
timestamp 1644511149
transform 1 0 39376 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_433
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_445
timestamp 1644511149
transform 1 0 42044 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_457
timestamp 1644511149
transform 1 0 43148 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_489
timestamp 1644511149
transform 1 0 46092 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_501
timestamp 1644511149
transform 1 0 47196 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_507
timestamp 1644511149
transform 1 0 47748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_512
timestamp 1644511149
transform 1 0 48208 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_43_6
timestamp 1644511149
transform 1 0 1656 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_27
timestamp 1644511149
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_39
timestamp 1644511149
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_51
timestamp 1644511149
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_55
timestamp 1644511149
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_43_64
timestamp 1644511149
transform 1 0 6992 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_68
timestamp 1644511149
transform 1 0 7360 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_76
timestamp 1644511149
transform 1 0 8096 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_80
timestamp 1644511149
transform 1 0 8464 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_88
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_99
timestamp 1644511149
transform 1 0 10212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_120
timestamp 1644511149
transform 1 0 12144 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_128
timestamp 1644511149
transform 1 0 12880 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_133
timestamp 1644511149
transform 1 0 13340 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_141
timestamp 1644511149
transform 1 0 14076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_145
timestamp 1644511149
transform 1 0 14444 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_157
timestamp 1644511149
transform 1 0 15548 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_165
timestamp 1644511149
transform 1 0 16284 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_175
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_183
timestamp 1644511149
transform 1 0 17940 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_202
timestamp 1644511149
transform 1 0 19688 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_212
timestamp 1644511149
transform 1 0 20608 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_237
timestamp 1644511149
transform 1 0 22908 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_249
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_253
timestamp 1644511149
transform 1 0 24380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_263
timestamp 1644511149
transform 1 0 25300 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_276
timestamp 1644511149
transform 1 0 26496 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_286
timestamp 1644511149
transform 1 0 27416 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_299
timestamp 1644511149
transform 1 0 28612 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_307
timestamp 1644511149
transform 1 0 29348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_329
timestamp 1644511149
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_335
timestamp 1644511149
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_341
timestamp 1644511149
transform 1 0 32476 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_366
timestamp 1644511149
transform 1 0 34776 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_382
timestamp 1644511149
transform 1 0 36248 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_390
timestamp 1644511149
transform 1 0 36984 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_393
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_405
timestamp 1644511149
transform 1 0 38364 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_417
timestamp 1644511149
transform 1 0 39468 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_429
timestamp 1644511149
transform 1 0 40572 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_441
timestamp 1644511149
transform 1 0 41676 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_447
timestamp 1644511149
transform 1 0 42228 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_461
timestamp 1644511149
transform 1 0 43516 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_473
timestamp 1644511149
transform 1 0 44620 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_485
timestamp 1644511149
transform 1 0 45724 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_497
timestamp 1644511149
transform 1 0 46828 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_503
timestamp 1644511149
transform 1 0 47380 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_43_505
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_513
timestamp 1644511149
transform 1 0 48300 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_44_24
timestamp 1644511149
transform 1 0 3312 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_29
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_41
timestamp 1644511149
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_53
timestamp 1644511149
transform 1 0 5980 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_80
timestamp 1644511149
transform 1 0 8464 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_106
timestamp 1644511149
transform 1 0 10856 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_118
timestamp 1644511149
transform 1 0 11960 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_130
timestamp 1644511149
transform 1 0 13064 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1644511149
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_141
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_149
timestamp 1644511149
transform 1 0 14812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_44_171
timestamp 1644511149
transform 1 0 16836 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_197
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_204
timestamp 1644511149
transform 1 0 19872 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_216
timestamp 1644511149
transform 1 0 20976 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_228
timestamp 1644511149
transform 1 0 22080 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_240
timestamp 1644511149
transform 1 0 23184 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_253
timestamp 1644511149
transform 1 0 24380 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_263
timestamp 1644511149
transform 1 0 25300 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_280
timestamp 1644511149
transform 1 0 26864 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_44_287
timestamp 1644511149
transform 1 0 27508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_44_292
timestamp 1644511149
transform 1 0 27968 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_304
timestamp 1644511149
transform 1 0 29072 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_313
timestamp 1644511149
transform 1 0 29900 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_326
timestamp 1644511149
transform 1 0 31096 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_346
timestamp 1644511149
transform 1 0 32936 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_350
timestamp 1644511149
transform 1 0 33304 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_369
timestamp 1644511149
transform 1 0 35052 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_373
timestamp 1644511149
transform 1 0 35420 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_395
timestamp 1644511149
transform 1 0 37444 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_407
timestamp 1644511149
transform 1 0 38548 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_419
timestamp 1644511149
transform 1 0 39652 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_433
timestamp 1644511149
transform 1 0 40940 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_445
timestamp 1644511149
transform 1 0 42044 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_457
timestamp 1644511149
transform 1 0 43148 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_469
timestamp 1644511149
transform 1 0 44252 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_507
timestamp 1644511149
transform 1 0 47748 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_512
timestamp 1644511149
transform 1 0 48208 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_28
timestamp 1644511149
transform 1 0 3680 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_40
timestamp 1644511149
transform 1 0 4784 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_68
timestamp 1644511149
transform 1 0 7360 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_45_81
timestamp 1644511149
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_93
timestamp 1644511149
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_105
timestamp 1644511149
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_111
timestamp 1644511149
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_125
timestamp 1644511149
transform 1 0 12604 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_140
timestamp 1644511149
transform 1 0 13984 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_150
timestamp 1644511149
transform 1 0 14904 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_156
timestamp 1644511149
transform 1 0 15456 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_163
timestamp 1644511149
transform 1 0 16100 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_167
timestamp 1644511149
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_173
timestamp 1644511149
transform 1 0 17020 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_178
timestamp 1644511149
transform 1 0 17480 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_45_190
timestamp 1644511149
transform 1 0 18584 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_198
timestamp 1644511149
transform 1 0 19320 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_207
timestamp 1644511149
transform 1 0 20148 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1644511149
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_45_254
timestamp 1644511149
transform 1 0 24472 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_276
timestamp 1644511149
transform 1 0 26496 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_297
timestamp 1644511149
transform 1 0 28428 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_301
timestamp 1644511149
transform 1 0 28796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_310
timestamp 1644511149
transform 1 0 29624 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_332
timestamp 1644511149
transform 1 0 31648 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_342
timestamp 1644511149
transform 1 0 32568 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_367
timestamp 1644511149
transform 1 0 34868 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_375
timestamp 1644511149
transform 1 0 35604 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_383
timestamp 1644511149
transform 1 0 36340 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_396
timestamp 1644511149
transform 1 0 37536 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_403
timestamp 1644511149
transform 1 0 38180 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_415
timestamp 1644511149
transform 1 0 39284 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_427
timestamp 1644511149
transform 1 0 40388 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_439
timestamp 1644511149
transform 1 0 41492 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_447
timestamp 1644511149
transform 1 0 42228 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_473
timestamp 1644511149
transform 1 0 44620 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_485
timestamp 1644511149
transform 1 0 45724 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_497
timestamp 1644511149
transform 1 0 46828 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_503
timestamp 1644511149
transform 1 0 47380 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_513
timestamp 1644511149
transform 1 0 48300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_6
timestamp 1644511149
transform 1 0 1656 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_13
timestamp 1644511149
transform 1 0 2300 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_20
timestamp 1644511149
transform 1 0 2944 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_61
timestamp 1644511149
transform 1 0 6716 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_78
timestamp 1644511149
transform 1 0 8280 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_93
timestamp 1644511149
transform 1 0 9660 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_97
timestamp 1644511149
transform 1 0 10028 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_101
timestamp 1644511149
transform 1 0 10396 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_110
timestamp 1644511149
transform 1 0 11224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_130
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_138
timestamp 1644511149
transform 1 0 13800 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_141
timestamp 1644511149
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_153
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_169
timestamp 1644511149
transform 1 0 16652 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_177
timestamp 1644511149
transform 1 0 17388 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_183
timestamp 1644511149
transform 1 0 17940 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_192
timestamp 1644511149
transform 1 0 18768 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_201
timestamp 1644511149
transform 1 0 19596 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_218
timestamp 1644511149
transform 1 0 21160 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_238
timestamp 1644511149
transform 1 0 23000 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1644511149
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_280
timestamp 1644511149
transform 1 0 26864 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_301
timestamp 1644511149
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_325
timestamp 1644511149
transform 1 0 31004 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_329
timestamp 1644511149
transform 1 0 31372 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_336
timestamp 1644511149
transform 1 0 32016 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_360
timestamp 1644511149
transform 1 0 34224 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_369
timestamp 1644511149
transform 1 0 35052 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_396
timestamp 1644511149
transform 1 0 37536 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1644511149
transform 1 0 38640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_445
timestamp 1644511149
transform 1 0 42044 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_457
timestamp 1644511149
transform 1 0 43148 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_469
timestamp 1644511149
transform 1 0 44252 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_475
timestamp 1644511149
transform 1 0 44804 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_477
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_489
timestamp 1644511149
transform 1 0 46092 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_501
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_513
timestamp 1644511149
transform 1 0 48300 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_15
timestamp 1644511149
transform 1 0 2484 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_38
timestamp 1644511149
transform 1 0 4600 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_50
timestamp 1644511149
transform 1 0 5704 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_47_89
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_108
timestamp 1644511149
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_123
timestamp 1644511149
transform 1 0 12420 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_127
timestamp 1644511149
transform 1 0 12788 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_131
timestamp 1644511149
transform 1 0 13156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_139
timestamp 1644511149
transform 1 0 13892 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_145
timestamp 1644511149
transform 1 0 14444 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_159
timestamp 1644511149
transform 1 0 15732 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_167
timestamp 1644511149
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_169
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_177
timestamp 1644511149
transform 1 0 17388 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_47_223
timestamp 1644511149
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_231
timestamp 1644511149
transform 1 0 22356 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_235
timestamp 1644511149
transform 1 0 22724 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_250
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_258
timestamp 1644511149
transform 1 0 24840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_270
timestamp 1644511149
transform 1 0 25944 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_278
timestamp 1644511149
transform 1 0 26680 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_301
timestamp 1644511149
transform 1 0 28796 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_311
timestamp 1644511149
transform 1 0 29716 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_319
timestamp 1644511149
transform 1 0 30452 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_332
timestamp 1644511149
transform 1 0 31648 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_47_359
timestamp 1644511149
transform 1 0 34132 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_384
timestamp 1644511149
transform 1 0 36432 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_396
timestamp 1644511149
transform 1 0 37536 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_408
timestamp 1644511149
transform 1 0 38640 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_420
timestamp 1644511149
transform 1 0 39744 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_432
timestamp 1644511149
transform 1 0 40848 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_444
timestamp 1644511149
transform 1 0 41952 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_449
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_461
timestamp 1644511149
transform 1 0 43516 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_485
timestamp 1644511149
transform 1 0 45724 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_497
timestamp 1644511149
transform 1 0 46828 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_503
timestamp 1644511149
transform 1 0 47380 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_47_512
timestamp 1644511149
transform 1 0 48208 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_24
timestamp 1644511149
transform 1 0 3312 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_65
timestamp 1644511149
transform 1 0 7084 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_73
timestamp 1644511149
transform 1 0 7820 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_80
timestamp 1644511149
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_93
timestamp 1644511149
transform 1 0 9660 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_101
timestamp 1644511149
transform 1 0 10396 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_112
timestamp 1644511149
transform 1 0 11408 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_125
timestamp 1644511149
transform 1 0 12604 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_132
timestamp 1644511149
transform 1 0 13248 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_48_148
timestamp 1644511149
transform 1 0 14720 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_156
timestamp 1644511149
transform 1 0 15456 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_169
timestamp 1644511149
transform 1 0 16652 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_179
timestamp 1644511149
transform 1 0 17572 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_183
timestamp 1644511149
transform 1 0 17940 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_48_197
timestamp 1644511149
transform 1 0 19228 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_215
timestamp 1644511149
transform 1 0 20884 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_227
timestamp 1644511149
transform 1 0 21988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_239
timestamp 1644511149
transform 1 0 23092 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_243
timestamp 1644511149
transform 1 0 23460 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_257
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_263
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_268
timestamp 1644511149
transform 1 0 25760 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_282
timestamp 1644511149
transform 1 0 27048 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_48_297
timestamp 1644511149
transform 1 0 28428 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_305
timestamp 1644511149
transform 1 0 29164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1644511149
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_48_343
timestamp 1644511149
transform 1 0 32660 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_358
timestamp 1644511149
transform 1 0 34040 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_48_368
timestamp 1644511149
transform 1 0 34960 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_48_395
timestamp 1644511149
transform 1 0 37444 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_407
timestamp 1644511149
transform 1 0 38548 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_445
timestamp 1644511149
transform 1 0 42044 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_457
timestamp 1644511149
transform 1 0 43148 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_469
timestamp 1644511149
transform 1 0 44252 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_48_489
timestamp 1644511149
transform 1 0 46092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_48_512
timestamp 1644511149
transform 1 0 48208 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_9
timestamp 1644511149
transform 1 0 1932 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_16
timestamp 1644511149
transform 1 0 2576 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_23
timestamp 1644511149
transform 1 0 3220 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_35
timestamp 1644511149
transform 1 0 4324 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_47
timestamp 1644511149
transform 1 0 5428 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_55
timestamp 1644511149
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_93
timestamp 1644511149
transform 1 0 9660 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_98
timestamp 1644511149
transform 1 0 10120 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_107
timestamp 1644511149
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_111
timestamp 1644511149
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_117
timestamp 1644511149
transform 1 0 11868 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_125
timestamp 1644511149
transform 1 0 12604 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_142
timestamp 1644511149
transform 1 0 14168 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_150
timestamp 1644511149
transform 1 0 14904 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_164
timestamp 1644511149
transform 1 0 16192 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_185
timestamp 1644511149
transform 1 0 18124 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_193
timestamp 1644511149
transform 1 0 18860 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_200
timestamp 1644511149
transform 1 0 19504 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_212
timestamp 1644511149
transform 1 0 20608 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_237
timestamp 1644511149
transform 1 0 22908 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_241
timestamp 1644511149
transform 1 0 23276 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_263
timestamp 1644511149
transform 1 0 25300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_270
timestamp 1644511149
transform 1 0 25944 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_278
timestamp 1644511149
transform 1 0 26680 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_49_281
timestamp 1644511149
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_293
timestamp 1644511149
transform 1 0 28060 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_49_315
timestamp 1644511149
transform 1 0 30084 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_49_331
timestamp 1644511149
transform 1 0 31556 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_354
timestamp 1644511149
transform 1 0 33672 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_362
timestamp 1644511149
transform 1 0 34408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_384
timestamp 1644511149
transform 1 0 36432 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_49_396
timestamp 1644511149
transform 1 0 37536 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_408
timestamp 1644511149
transform 1 0 38640 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_420
timestamp 1644511149
transform 1 0 39744 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_432
timestamp 1644511149
transform 1 0 40848 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_444
timestamp 1644511149
transform 1 0 41952 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_461
timestamp 1644511149
transform 1 0 43516 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_473
timestamp 1644511149
transform 1 0 44620 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_485
timestamp 1644511149
transform 1 0 45724 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_500
timestamp 1644511149
transform 1 0 47104 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_508
timestamp 1644511149
transform 1 0 47840 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_50_24
timestamp 1644511149
transform 1 0 3312 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_29
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_41
timestamp 1644511149
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_53
timestamp 1644511149
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_65
timestamp 1644511149
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_77
timestamp 1644511149
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_83
timestamp 1644511149
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_96
timestamp 1644511149
transform 1 0 9936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_109
timestamp 1644511149
transform 1 0 11132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_123
timestamp 1644511149
transform 1 0 12420 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_135
timestamp 1644511149
transform 1 0 13524 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_139
timestamp 1644511149
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_156
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_187
timestamp 1644511149
transform 1 0 18308 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_50_195
timestamp 1644511149
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_197
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_205
timestamp 1644511149
transform 1 0 19964 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_229
timestamp 1644511149
transform 1 0 22172 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_241
timestamp 1644511149
transform 1 0 23276 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_249
timestamp 1644511149
transform 1 0 24012 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_253
timestamp 1644511149
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_265
timestamp 1644511149
transform 1 0 25484 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_284
timestamp 1644511149
transform 1 0 27232 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_297
timestamp 1644511149
transform 1 0 28428 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_50_305
timestamp 1644511149
transform 1 0 29164 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_329
timestamp 1644511149
transform 1 0 31372 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_349
timestamp 1644511149
transform 1 0 33212 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_356
timestamp 1644511149
transform 1 0 33856 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_50_368
timestamp 1644511149
transform 1 0 34960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_395
timestamp 1644511149
transform 1 0 37444 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_407
timestamp 1644511149
transform 1 0 38548 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_419
timestamp 1644511149
transform 1 0 39652 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_457
timestamp 1644511149
transform 1 0 43148 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_469
timestamp 1644511149
transform 1 0 44252 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_475
timestamp 1644511149
transform 1 0 44804 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_477
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_489
timestamp 1644511149
transform 1 0 46092 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_501
timestamp 1644511149
transform 1 0 47196 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_512
timestamp 1644511149
transform 1 0 48208 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_8
timestamp 1644511149
transform 1 0 1840 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_69
timestamp 1644511149
transform 1 0 7452 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_88
timestamp 1644511149
transform 1 0 9200 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_108
timestamp 1644511149
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_124
timestamp 1644511149
transform 1 0 12512 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_51_139
timestamp 1644511149
transform 1 0 13892 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_149
timestamp 1644511149
transform 1 0 14812 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_157
timestamp 1644511149
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_165
timestamp 1644511149
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_173
timestamp 1644511149
transform 1 0 17020 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_177
timestamp 1644511149
transform 1 0 17388 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_181
timestamp 1644511149
transform 1 0 17756 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_204
timestamp 1644511149
transform 1 0 19872 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_212
timestamp 1644511149
transform 1 0 20608 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_220
timestamp 1644511149
transform 1 0 21344 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_253
timestamp 1644511149
transform 1 0 24380 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_270
timestamp 1644511149
transform 1 0 25944 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_278
timestamp 1644511149
transform 1 0 26680 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_293
timestamp 1644511149
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_305
timestamp 1644511149
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_317
timestamp 1644511149
transform 1 0 30268 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_323
timestamp 1644511149
transform 1 0 30820 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_342
timestamp 1644511149
transform 1 0 32568 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_350
timestamp 1644511149
transform 1 0 33304 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_372
timestamp 1644511149
transform 1 0 35328 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_384
timestamp 1644511149
transform 1 0 36432 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_393
timestamp 1644511149
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_405
timestamp 1644511149
transform 1 0 38364 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_417
timestamp 1644511149
transform 1 0 39468 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_429
timestamp 1644511149
transform 1 0 40572 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_441
timestamp 1644511149
transform 1 0 41676 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_449
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_461
timestamp 1644511149
transform 1 0 43516 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_473
timestamp 1644511149
transform 1 0 44620 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_485
timestamp 1644511149
transform 1 0 45724 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_497
timestamp 1644511149
transform 1 0 46828 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_51_513
timestamp 1644511149
transform 1 0 48300 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_11
timestamp 1644511149
transform 1 0 2116 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_22
timestamp 1644511149
transform 1 0 3128 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_77
timestamp 1644511149
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_83
timestamp 1644511149
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_97
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_102
timestamp 1644511149
transform 1 0 10488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_114
timestamp 1644511149
transform 1 0 11592 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_126
timestamp 1644511149
transform 1 0 12696 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_138
timestamp 1644511149
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_52_146
timestamp 1644511149
transform 1 0 14536 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_154
timestamp 1644511149
transform 1 0 15272 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_166
timestamp 1644511149
transform 1 0 16376 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_175
timestamp 1644511149
transform 1 0 17204 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_182
timestamp 1644511149
transform 1 0 17848 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_194
timestamp 1644511149
transform 1 0 18952 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_201
timestamp 1644511149
transform 1 0 19596 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_52_232
timestamp 1644511149
transform 1 0 22448 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_244
timestamp 1644511149
transform 1 0 23552 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_262
timestamp 1644511149
transform 1 0 25208 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_274
timestamp 1644511149
transform 1 0 26312 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_280
timestamp 1644511149
transform 1 0 26864 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_297
timestamp 1644511149
transform 1 0 28428 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_305
timestamp 1644511149
transform 1 0 29164 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_334
timestamp 1644511149
transform 1 0 31832 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_346
timestamp 1644511149
transform 1 0 32936 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_352
timestamp 1644511149
transform 1 0 33488 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_356
timestamp 1644511149
transform 1 0 33856 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_360
timestamp 1644511149
transform 1 0 34224 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_386
timestamp 1644511149
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_398
timestamp 1644511149
transform 1 0 37720 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_410
timestamp 1644511149
transform 1 0 38824 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_418
timestamp 1644511149
transform 1 0 39560 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_52_429
timestamp 1644511149
transform 1 0 40572 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_435
timestamp 1644511149
transform 1 0 41124 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_447
timestamp 1644511149
transform 1 0 42228 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_459
timestamp 1644511149
transform 1 0 43332 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_471
timestamp 1644511149
transform 1 0 44436 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_477
timestamp 1644511149
transform 1 0 44988 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_489
timestamp 1644511149
transform 1 0 46092 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_501
timestamp 1644511149
transform 1 0 47196 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_513
timestamp 1644511149
transform 1 0 48300 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_32
timestamp 1644511149
transform 1 0 4048 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_44
timestamp 1644511149
transform 1 0 5152 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_69
timestamp 1644511149
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_81
timestamp 1644511149
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_105
timestamp 1644511149
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_129
timestamp 1644511149
transform 1 0 12972 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_139
timestamp 1644511149
transform 1 0 13892 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_148
timestamp 1644511149
transform 1 0 14720 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_160
timestamp 1644511149
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_185
timestamp 1644511149
transform 1 0 18124 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_197
timestamp 1644511149
transform 1 0 19228 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_205
timestamp 1644511149
transform 1 0 19964 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_214
timestamp 1644511149
transform 1 0 20792 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_222
timestamp 1644511149
transform 1 0 21528 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_53_225
timestamp 1644511149
transform 1 0 21804 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_231
timestamp 1644511149
transform 1 0 22356 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_237
timestamp 1644511149
transform 1 0 22908 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_243
timestamp 1644511149
transform 1 0 23460 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_249
timestamp 1644511149
transform 1 0 24012 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_254
timestamp 1644511149
transform 1 0 24472 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_264
timestamp 1644511149
transform 1 0 25392 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_272
timestamp 1644511149
transform 1 0 26128 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_285
timestamp 1644511149
transform 1 0 27324 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_297
timestamp 1644511149
transform 1 0 28428 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_307
timestamp 1644511149
transform 1 0 29348 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_319
timestamp 1644511149
transform 1 0 30452 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_331
timestamp 1644511149
transform 1 0 31556 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_335
timestamp 1644511149
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_345
timestamp 1644511149
transform 1 0 32844 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_357
timestamp 1644511149
transform 1 0 33948 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_369
timestamp 1644511149
transform 1 0 35052 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_381
timestamp 1644511149
transform 1 0 36156 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_53_389
timestamp 1644511149
transform 1 0 36892 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_393
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_405
timestamp 1644511149
transform 1 0 38364 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_417
timestamp 1644511149
transform 1 0 39468 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_429
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_441
timestamp 1644511149
transform 1 0 41676 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_447
timestamp 1644511149
transform 1 0 42228 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_473
timestamp 1644511149
transform 1 0 44620 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_485
timestamp 1644511149
transform 1 0 45724 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_497
timestamp 1644511149
transform 1 0 46828 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_503
timestamp 1644511149
transform 1 0 47380 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_53_512
timestamp 1644511149
transform 1 0 48208 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_32
timestamp 1644511149
transform 1 0 4048 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_44
timestamp 1644511149
transform 1 0 5152 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_56
timestamp 1644511149
transform 1 0 6256 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_68
timestamp 1644511149
transform 1 0 7360 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_85
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_93
timestamp 1644511149
transform 1 0 9660 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_102
timestamp 1644511149
transform 1 0 10488 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_114
timestamp 1644511149
transform 1 0 11592 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_151
timestamp 1644511149
transform 1 0 14996 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_163
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_171
timestamp 1644511149
transform 1 0 16836 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_176
timestamp 1644511149
transform 1 0 17296 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_185
timestamp 1644511149
transform 1 0 18124 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_193
timestamp 1644511149
transform 1 0 18860 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_222
timestamp 1644511149
transform 1 0 21528 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_234
timestamp 1644511149
transform 1 0 22632 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_246
timestamp 1644511149
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_253
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_265
timestamp 1644511149
transform 1 0 25484 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_271
timestamp 1644511149
transform 1 0 26036 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_280
timestamp 1644511149
transform 1 0 26864 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_289
timestamp 1644511149
transform 1 0 27692 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_302
timestamp 1644511149
transform 1 0 28888 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_54_314
timestamp 1644511149
transform 1 0 29992 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_54_334
timestamp 1644511149
transform 1 0 31832 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_340
timestamp 1644511149
transform 1 0 32384 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_357
timestamp 1644511149
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_363
timestamp 1644511149
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_54_365
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_374
timestamp 1644511149
transform 1 0 35512 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_386
timestamp 1644511149
transform 1 0 36616 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_410
timestamp 1644511149
transform 1 0 38824 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_418
timestamp 1644511149
transform 1 0 39560 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_445
timestamp 1644511149
transform 1 0 42044 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_457
timestamp 1644511149
transform 1 0 43148 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_469
timestamp 1644511149
transform 1 0 44252 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_475
timestamp 1644511149
transform 1 0 44804 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_489
timestamp 1644511149
transform 1 0 46092 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_501
timestamp 1644511149
transform 1 0 47196 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_512
timestamp 1644511149
transform 1 0 48208 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_28
timestamp 1644511149
transform 1 0 3680 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_40
timestamp 1644511149
transform 1 0 4784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_52
timestamp 1644511149
transform 1 0 5888 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_69
timestamp 1644511149
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_81
timestamp 1644511149
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_130
timestamp 1644511149
transform 1 0 13064 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_134
timestamp 1644511149
transform 1 0 13432 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_138
timestamp 1644511149
transform 1 0 13800 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_159
timestamp 1644511149
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_167
timestamp 1644511149
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_177
timestamp 1644511149
transform 1 0 17388 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_186
timestamp 1644511149
transform 1 0 18216 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_55_198
timestamp 1644511149
transform 1 0 19320 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_217
timestamp 1644511149
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_223
timestamp 1644511149
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_241
timestamp 1644511149
transform 1 0 23276 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_247
timestamp 1644511149
transform 1 0 23828 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_264
timestamp 1644511149
transform 1 0 25392 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_275
timestamp 1644511149
transform 1 0 26404 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_279
timestamp 1644511149
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_55_281
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 1644511149
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_55_292
timestamp 1644511149
transform 1 0 27968 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_301
timestamp 1644511149
transform 1 0 28796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_314
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1644511149
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_343
timestamp 1644511149
transform 1 0 32660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_355
timestamp 1644511149
transform 1 0 33764 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_367
timestamp 1644511149
transform 1 0 34868 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_379
timestamp 1644511149
transform 1 0 35972 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_55_391
timestamp 1644511149
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_393
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_405
timestamp 1644511149
transform 1 0 38364 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_417
timestamp 1644511149
transform 1 0 39468 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_429
timestamp 1644511149
transform 1 0 40572 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_441
timestamp 1644511149
transform 1 0 41676 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_447
timestamp 1644511149
transform 1 0 42228 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_461
timestamp 1644511149
transform 1 0 43516 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_473
timestamp 1644511149
transform 1 0 44620 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_513
timestamp 1644511149
transform 1 0 48300 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_11
timestamp 1644511149
transform 1 0 2116 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_23
timestamp 1644511149
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_65
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_77
timestamp 1644511149
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_83
timestamp 1644511149
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_85
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_97
timestamp 1644511149
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_109
timestamp 1644511149
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_121
timestamp 1644511149
transform 1 0 12236 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_136
timestamp 1644511149
transform 1 0 13616 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_149
timestamp 1644511149
transform 1 0 14812 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_161
timestamp 1644511149
transform 1 0 15916 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_165
timestamp 1644511149
transform 1 0 16284 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_182
timestamp 1644511149
transform 1 0 17848 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_192
timestamp 1644511149
transform 1 0 18768 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_197
timestamp 1644511149
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_209
timestamp 1644511149
transform 1 0 20332 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_222
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_239
timestamp 1644511149
transform 1 0 23092 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_248
timestamp 1644511149
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_56_262
timestamp 1644511149
transform 1 0 25208 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_284
timestamp 1644511149
transform 1 0 27232 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_292
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_304
timestamp 1644511149
transform 1 0 29072 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_318
timestamp 1644511149
transform 1 0 30360 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_330
timestamp 1644511149
transform 1 0 31464 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_343
timestamp 1644511149
transform 1 0 32660 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_355
timestamp 1644511149
transform 1 0 33764 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_363
timestamp 1644511149
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_365
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_369
timestamp 1644511149
transform 1 0 35052 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_391
timestamp 1644511149
transform 1 0 37076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_403
timestamp 1644511149
transform 1 0 38180 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_415
timestamp 1644511149
transform 1 0 39284 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_419
timestamp 1644511149
transform 1 0 39652 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_477
timestamp 1644511149
transform 1 0 44988 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_489
timestamp 1644511149
transform 1 0 46092 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_56_512
timestamp 1644511149
transform 1 0 48208 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_9
timestamp 1644511149
transform 1 0 1932 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_13
timestamp 1644511149
transform 1 0 2300 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_20
timestamp 1644511149
transform 1 0 2944 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_32
timestamp 1644511149
transform 1 0 4048 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_44
timestamp 1644511149
transform 1 0 5152 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_69
timestamp 1644511149
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_81
timestamp 1644511149
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_93
timestamp 1644511149
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_105
timestamp 1644511149
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_111
timestamp 1644511149
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_125
timestamp 1644511149
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_137
timestamp 1644511149
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_149
timestamp 1644511149
transform 1 0 14812 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_155
timestamp 1644511149
transform 1 0 15364 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_164
timestamp 1644511149
transform 1 0 16192 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_173
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_176
timestamp 1644511149
transform 1 0 17296 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_183
timestamp 1644511149
transform 1 0 17940 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_191
timestamp 1644511149
transform 1 0 18676 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_199
timestamp 1644511149
transform 1 0 19412 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_205
timestamp 1644511149
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_217
timestamp 1644511149
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_223
timestamp 1644511149
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_241
timestamp 1644511149
transform 1 0 23276 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_57_250
timestamp 1644511149
transform 1 0 24104 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_258
timestamp 1644511149
transform 1 0 24840 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_269
timestamp 1644511149
transform 1 0 25852 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_277
timestamp 1644511149
transform 1 0 26588 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_281
timestamp 1644511149
transform 1 0 26956 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_289
timestamp 1644511149
transform 1 0 27692 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_295
timestamp 1644511149
transform 1 0 28244 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_308
timestamp 1644511149
transform 1 0 29440 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_314
timestamp 1644511149
transform 1 0 29992 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_331
timestamp 1644511149
transform 1 0 31556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_335
timestamp 1644511149
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_345
timestamp 1644511149
transform 1 0 32844 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_353
timestamp 1644511149
transform 1 0 33580 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_365
timestamp 1644511149
transform 1 0 34684 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_377
timestamp 1644511149
transform 1 0 35788 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_389
timestamp 1644511149
transform 1 0 36892 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_449
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_461
timestamp 1644511149
transform 1 0 43516 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_473
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_490
timestamp 1644511149
transform 1 0 46184 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_512
timestamp 1644511149
transform 1 0 48208 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_24
timestamp 1644511149
transform 1 0 3312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_77
timestamp 1644511149
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_83
timestamp 1644511149
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_97
timestamp 1644511149
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_121
timestamp 1644511149
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_133
timestamp 1644511149
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_139
timestamp 1644511149
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_58_149
timestamp 1644511149
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_58_166
timestamp 1644511149
transform 1 0 16376 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_174
timestamp 1644511149
transform 1 0 17112 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_186
timestamp 1644511149
transform 1 0 18216 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_197
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_209
timestamp 1644511149
transform 1 0 20332 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_217
timestamp 1644511149
transform 1 0 21068 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_230
timestamp 1644511149
transform 1 0 22264 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_242
timestamp 1644511149
transform 1 0 23368 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_248
timestamp 1644511149
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_263
timestamp 1644511149
transform 1 0 25300 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_282
timestamp 1644511149
transform 1 0 27048 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_289
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_297
timestamp 1644511149
transform 1 0 28428 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_304
timestamp 1644511149
transform 1 0 29072 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_337
timestamp 1644511149
transform 1 0 32108 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_357
timestamp 1644511149
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_363
timestamp 1644511149
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_368
timestamp 1644511149
transform 1 0 34960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_380
timestamp 1644511149
transform 1 0 36064 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_392
timestamp 1644511149
transform 1 0 37168 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_404
timestamp 1644511149
transform 1 0 38272 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_416
timestamp 1644511149
transform 1 0 39376 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_433
timestamp 1644511149
transform 1 0 40940 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_445
timestamp 1644511149
transform 1 0 42044 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_457
timestamp 1644511149
transform 1 0 43148 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_477
timestamp 1644511149
transform 1 0 44988 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_489
timestamp 1644511149
transform 1 0 46092 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_512
timestamp 1644511149
transform 1 0 48208 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_7
timestamp 1644511149
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_11
timestamp 1644511149
transform 1 0 2116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_23
timestamp 1644511149
transform 1 0 3220 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_35
timestamp 1644511149
transform 1 0 4324 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_47
timestamp 1644511149
transform 1 0 5428 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_69
timestamp 1644511149
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_81
timestamp 1644511149
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_93
timestamp 1644511149
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_105
timestamp 1644511149
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_111
timestamp 1644511149
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_116
timestamp 1644511149
transform 1 0 11776 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_128
timestamp 1644511149
transform 1 0 12880 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_140
timestamp 1644511149
transform 1 0 13984 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_152
timestamp 1644511149
transform 1 0 15088 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_169
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_197
timestamp 1644511149
transform 1 0 19228 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_204
timestamp 1644511149
transform 1 0 19872 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_220
timestamp 1644511149
transform 1 0 21344 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_241
timestamp 1644511149
transform 1 0 23276 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_255
timestamp 1644511149
transform 1 0 24564 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_268
timestamp 1644511149
transform 1 0 25760 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_276
timestamp 1644511149
transform 1 0 26496 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_285
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_300
timestamp 1644511149
transform 1 0 28704 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_312
timestamp 1644511149
transform 1 0 29808 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_324
timestamp 1644511149
transform 1 0 30912 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_332
timestamp 1644511149
transform 1 0 31648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_353
timestamp 1644511149
transform 1 0 33580 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_59_382
timestamp 1644511149
transform 1 0 36248 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_390
timestamp 1644511149
transform 1 0 36984 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_405
timestamp 1644511149
transform 1 0 38364 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_417
timestamp 1644511149
transform 1 0 39468 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_429
timestamp 1644511149
transform 1 0 40572 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_59_441
timestamp 1644511149
transform 1 0 41676 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_59_447
timestamp 1644511149
transform 1 0 42228 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_461
timestamp 1644511149
transform 1 0 43516 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_473
timestamp 1644511149
transform 1 0 44620 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_485
timestamp 1644511149
transform 1 0 45724 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_489
timestamp 1644511149
transform 1 0 46092 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_493
timestamp 1644511149
transform 1 0 46460 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_500
timestamp 1644511149
transform 1 0 47104 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_508
timestamp 1644511149
transform 1 0 47840 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_13
timestamp 1644511149
transform 1 0 2300 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_25
timestamp 1644511149
transform 1 0 3404 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_65
timestamp 1644511149
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_77
timestamp 1644511149
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_83
timestamp 1644511149
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_85
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_97
timestamp 1644511149
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_109
timestamp 1644511149
transform 1 0 11132 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_60_159
timestamp 1644511149
transform 1 0 15732 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_171
timestamp 1644511149
transform 1 0 16836 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_60_179
timestamp 1644511149
transform 1 0 17572 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_60_188
timestamp 1644511149
transform 1 0 18400 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_206
timestamp 1644511149
transform 1 0 20056 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_215
timestamp 1644511149
transform 1 0 20884 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_227
timestamp 1644511149
transform 1 0 21988 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_60_250
timestamp 1644511149
transform 1 0 24104 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_259
timestamp 1644511149
transform 1 0 24932 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_268
timestamp 1644511149
transform 1 0 25760 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_276
timestamp 1644511149
transform 1 0 26496 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_60_287
timestamp 1644511149
transform 1 0 27508 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_295
timestamp 1644511149
transform 1 0 28244 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_307
timestamp 1644511149
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_360
timestamp 1644511149
transform 1 0 34224 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_365
timestamp 1644511149
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_377
timestamp 1644511149
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_389
timestamp 1644511149
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_401
timestamp 1644511149
transform 1 0 37996 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_413
timestamp 1644511149
transform 1 0 39100 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_419
timestamp 1644511149
transform 1 0 39652 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_457
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_469
timestamp 1644511149
transform 1 0 44252 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_475
timestamp 1644511149
transform 1 0 44804 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_512
timestamp 1644511149
transform 1 0 48208 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_9
timestamp 1644511149
transform 1 0 1932 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_31
timestamp 1644511149
transform 1 0 3956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_43
timestamp 1644511149
transform 1 0 5060 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_57
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_69
timestamp 1644511149
transform 1 0 7452 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_74
timestamp 1644511149
transform 1 0 7912 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_86
timestamp 1644511149
transform 1 0 9016 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1644511149
transform 1 0 10120 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1644511149
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_125
timestamp 1644511149
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_137
timestamp 1644511149
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_149
timestamp 1644511149
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_161
timestamp 1644511149
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_167
timestamp 1644511149
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_173
timestamp 1644511149
transform 1 0 17020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_178
timestamp 1644511149
transform 1 0 17480 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_198
timestamp 1644511149
transform 1 0 19320 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_210
timestamp 1644511149
transform 1 0 20424 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_220
timestamp 1644511149
transform 1 0 21344 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_61_241
timestamp 1644511149
transform 1 0 23276 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_61_251
timestamp 1644511149
transform 1 0 24196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_61_262
timestamp 1644511149
transform 1 0 25208 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_275
timestamp 1644511149
transform 1 0 26404 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_301
timestamp 1644511149
transform 1 0 28796 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_313
timestamp 1644511149
transform 1 0 29900 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_325
timestamp 1644511149
transform 1 0 31004 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_61_333
timestamp 1644511149
transform 1 0 31740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_349
timestamp 1644511149
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_361
timestamp 1644511149
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_373
timestamp 1644511149
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_385
timestamp 1644511149
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_391
timestamp 1644511149
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_429
timestamp 1644511149
transform 1 0 40572 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_441
timestamp 1644511149
transform 1 0 41676 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_485
timestamp 1644511149
transform 1 0 45724 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_497
timestamp 1644511149
transform 1 0 46828 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_503
timestamp 1644511149
transform 1 0 47380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_508
timestamp 1644511149
transform 1 0 47840 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_3
timestamp 1644511149
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_15
timestamp 1644511149
transform 1 0 2484 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_23
timestamp 1644511149
transform 1 0 3220 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_61
timestamp 1644511149
transform 1 0 6716 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_62_78
timestamp 1644511149
transform 1 0 8280 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_62_85
timestamp 1644511149
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_97
timestamp 1644511149
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_109
timestamp 1644511149
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_121
timestamp 1644511149
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_133
timestamp 1644511149
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_139
timestamp 1644511149
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_171
timestamp 1644511149
transform 1 0 16836 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_176
timestamp 1644511149
transform 1 0 17296 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_188
timestamp 1644511149
transform 1 0 18400 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_202
timestamp 1644511149
transform 1 0 19688 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_206
timestamp 1644511149
transform 1 0 20056 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_210
timestamp 1644511149
transform 1 0 20424 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_219
timestamp 1644511149
transform 1 0 21252 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_232
timestamp 1644511149
transform 1 0 22448 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_240
timestamp 1644511149
transform 1 0 23184 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_247
timestamp 1644511149
transform 1 0 23828 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_251
timestamp 1644511149
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_62_253
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_62_260
timestamp 1644511149
transform 1 0 25024 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_268
timestamp 1644511149
transform 1 0 25760 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_275
timestamp 1644511149
transform 1 0 26404 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_279
timestamp 1644511149
transform 1 0 26772 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_309
timestamp 1644511149
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_321
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_333
timestamp 1644511149
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_357
timestamp 1644511149
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_363
timestamp 1644511149
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_377
timestamp 1644511149
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_389
timestamp 1644511149
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_401
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_413
timestamp 1644511149
transform 1 0 39100 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_419
timestamp 1644511149
transform 1 0 39652 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_421
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_433
timestamp 1644511149
transform 1 0 40940 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_445
timestamp 1644511149
transform 1 0 42044 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_457
timestamp 1644511149
transform 1 0 43148 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_469
timestamp 1644511149
transform 1 0 44252 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_475
timestamp 1644511149
transform 1 0 44804 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_489
timestamp 1644511149
transform 1 0 46092 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_501
timestamp 1644511149
transform 1 0 47196 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_507
timestamp 1644511149
transform 1 0 47748 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_512
timestamp 1644511149
transform 1 0 48208 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_3
timestamp 1644511149
transform 1 0 1380 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_14
timestamp 1644511149
transform 1 0 2392 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_26
timestamp 1644511149
transform 1 0 3496 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_38
timestamp 1644511149
transform 1 0 4600 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_50
timestamp 1644511149
transform 1 0 5704 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_63_57
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_65
timestamp 1644511149
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_87
timestamp 1644511149
transform 1 0 9108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_99
timestamp 1644511149
transform 1 0 10212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_111
timestamp 1644511149
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_149
timestamp 1644511149
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_161
timestamp 1644511149
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_189
timestamp 1644511149
transform 1 0 18492 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_206
timestamp 1644511149
transform 1 0 20056 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_214
timestamp 1644511149
transform 1 0 20792 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_222
timestamp 1644511149
transform 1 0 21528 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_63_252
timestamp 1644511149
transform 1 0 24288 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_63_272
timestamp 1644511149
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_63_285
timestamp 1644511149
transform 1 0 27324 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_289
timestamp 1644511149
transform 1 0 27692 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_306
timestamp 1644511149
transform 1 0 29256 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_316
timestamp 1644511149
transform 1 0 30176 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_328
timestamp 1644511149
transform 1 0 31280 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_63_337
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_349
timestamp 1644511149
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_361
timestamp 1644511149
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_373
timestamp 1644511149
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_385
timestamp 1644511149
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_391
timestamp 1644511149
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_405
timestamp 1644511149
transform 1 0 38364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_417
timestamp 1644511149
transform 1 0 39468 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_429
timestamp 1644511149
transform 1 0 40572 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_441
timestamp 1644511149
transform 1 0 41676 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_447
timestamp 1644511149
transform 1 0 42228 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_461
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_473
timestamp 1644511149
transform 1 0 44620 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_485
timestamp 1644511149
transform 1 0 45724 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1644511149
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_508
timestamp 1644511149
transform 1 0 47840 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_64_13
timestamp 1644511149
transform 1 0 2300 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_25
timestamp 1644511149
transform 1 0 3404 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_41
timestamp 1644511149
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_53
timestamp 1644511149
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_65
timestamp 1644511149
transform 1 0 7084 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_70
timestamp 1644511149
transform 1 0 7544 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_82
timestamp 1644511149
transform 1 0 8648 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_97
timestamp 1644511149
transform 1 0 10028 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_109
timestamp 1644511149
transform 1 0 11132 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_121
timestamp 1644511149
transform 1 0 12236 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_133
timestamp 1644511149
transform 1 0 13340 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_139
timestamp 1644511149
transform 1 0 13892 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_64_165
timestamp 1644511149
transform 1 0 16284 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_192
timestamp 1644511149
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_206
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_214
timestamp 1644511149
transform 1 0 20792 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_232
timestamp 1644511149
transform 1 0 22448 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_240
timestamp 1644511149
transform 1 0 23184 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_262
timestamp 1644511149
transform 1 0 25208 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_274
timestamp 1644511149
transform 1 0 26312 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_286
timestamp 1644511149
transform 1 0 27416 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_64_292
timestamp 1644511149
transform 1 0 27968 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_304
timestamp 1644511149
transform 1 0 29072 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_325
timestamp 1644511149
transform 1 0 31004 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_349
timestamp 1644511149
transform 1 0 33212 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_64_361
timestamp 1644511149
transform 1 0 34316 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_377
timestamp 1644511149
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_389
timestamp 1644511149
transform 1 0 36892 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_401
timestamp 1644511149
transform 1 0 37996 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_413
timestamp 1644511149
transform 1 0 39100 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_421
timestamp 1644511149
transform 1 0 39836 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_445
timestamp 1644511149
transform 1 0 42044 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_64_457
timestamp 1644511149
transform 1 0 43148 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_469
timestamp 1644511149
transform 1 0 44252 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_475
timestamp 1644511149
transform 1 0 44804 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_512
timestamp 1644511149
transform 1 0 48208 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_3
timestamp 1644511149
transform 1 0 1380 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_11
timestamp 1644511149
transform 1 0 2116 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_19
timestamp 1644511149
transform 1 0 2852 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_23
timestamp 1644511149
transform 1 0 3220 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_35
timestamp 1644511149
transform 1 0 4324 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_47
timestamp 1644511149
transform 1 0 5428 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_55
timestamp 1644511149
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_57
timestamp 1644511149
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_69
timestamp 1644511149
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_81
timestamp 1644511149
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_93
timestamp 1644511149
transform 1 0 9660 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_105
timestamp 1644511149
transform 1 0 10764 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_111
timestamp 1644511149
transform 1 0 11316 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_113
timestamp 1644511149
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_125
timestamp 1644511149
transform 1 0 12604 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_137
timestamp 1644511149
transform 1 0 13708 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_149
timestamp 1644511149
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_161
timestamp 1644511149
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_167
timestamp 1644511149
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_169
timestamp 1644511149
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_181
timestamp 1644511149
transform 1 0 17756 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_65_185
timestamp 1644511149
transform 1 0 18124 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_191
timestamp 1644511149
transform 1 0 18676 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_203
timestamp 1644511149
transform 1 0 19780 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_211
timestamp 1644511149
transform 1 0 20516 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_220
timestamp 1644511149
transform 1 0 21344 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_65_225
timestamp 1644511149
transform 1 0 21804 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_231
timestamp 1644511149
transform 1 0 22356 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_65_248
timestamp 1644511149
transform 1 0 23920 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_65_261
timestamp 1644511149
transform 1 0 25116 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_65_271
timestamp 1644511149
transform 1 0 26036 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_279
timestamp 1644511149
transform 1 0 26772 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_281
timestamp 1644511149
transform 1 0 26956 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_65_293
timestamp 1644511149
transform 1 0 28060 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_65_301
timestamp 1644511149
transform 1 0 28796 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_310
timestamp 1644511149
transform 1 0 29624 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_322
timestamp 1644511149
transform 1 0 30728 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_65_334
timestamp 1644511149
transform 1 0 31832 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_65_337
timestamp 1644511149
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_349
timestamp 1644511149
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_361
timestamp 1644511149
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_373
timestamp 1644511149
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_385
timestamp 1644511149
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_391
timestamp 1644511149
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_393
timestamp 1644511149
transform 1 0 37260 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_405
timestamp 1644511149
transform 1 0 38364 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_417
timestamp 1644511149
transform 1 0 39468 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_429
timestamp 1644511149
transform 1 0 40572 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_65_441
timestamp 1644511149
transform 1 0 41676 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_65_447
timestamp 1644511149
transform 1 0 42228 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_65_449
timestamp 1644511149
transform 1 0 42412 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_461
timestamp 1644511149
transform 1 0 43516 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_473
timestamp 1644511149
transform 1 0 44620 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_65_485
timestamp 1644511149
transform 1 0 45724 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_65_500
timestamp 1644511149
transform 1 0 47104 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_65_505
timestamp 1644511149
transform 1 0 47564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_65_512
timestamp 1644511149
transform 1 0 48208 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_66_3
timestamp 1644511149
transform 1 0 1380 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_66_14
timestamp 1644511149
transform 1 0 2392 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_26
timestamp 1644511149
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_66_29
timestamp 1644511149
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_41
timestamp 1644511149
transform 1 0 4876 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_53
timestamp 1644511149
transform 1 0 5980 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_65
timestamp 1644511149
transform 1 0 7084 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_77
timestamp 1644511149
transform 1 0 8188 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_83
timestamp 1644511149
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_85
timestamp 1644511149
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_97
timestamp 1644511149
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_109
timestamp 1644511149
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_121
timestamp 1644511149
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_133
timestamp 1644511149
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_139
timestamp 1644511149
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_141
timestamp 1644511149
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_153
timestamp 1644511149
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_165
timestamp 1644511149
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_66_177
timestamp 1644511149
transform 1 0 17388 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_66_182
timestamp 1644511149
transform 1 0 17848 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_190
timestamp 1644511149
transform 1 0 18584 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_66_197
timestamp 1644511149
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_205
timestamp 1644511149
transform 1 0 19964 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_217
timestamp 1644511149
transform 1 0 21068 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_66_225
timestamp 1644511149
transform 1 0 21804 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_235
timestamp 1644511149
transform 1 0 22724 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_66_245
timestamp 1644511149
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_251
timestamp 1644511149
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_66_253
timestamp 1644511149
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_66_264
timestamp 1644511149
transform 1 0 25392 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_66_276
timestamp 1644511149
transform 1 0 26496 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_66_284
timestamp 1644511149
transform 1 0 27232 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_66_292
timestamp 1644511149
transform 1 0 27968 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_66_304
timestamp 1644511149
transform 1 0 29072 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_66_325
timestamp 1644511149
transform 1 0 31004 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_337
timestamp 1644511149
transform 1 0 32108 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_349
timestamp 1644511149
transform 1 0 33212 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_66_361
timestamp 1644511149
transform 1 0 34316 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_66_365
timestamp 1644511149
transform 1 0 34684 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_377
timestamp 1644511149
transform 1 0 35788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_389
timestamp 1644511149
transform 1 0 36892 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_401
timestamp 1644511149
transform 1 0 37996 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_413
timestamp 1644511149
transform 1 0 39100 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_419
timestamp 1644511149
transform 1 0 39652 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_421
timestamp 1644511149
transform 1 0 39836 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_433
timestamp 1644511149
transform 1 0 40940 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_445
timestamp 1644511149
transform 1 0 42044 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_66_457
timestamp 1644511149
transform 1 0 43148 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_66_469
timestamp 1644511149
transform 1 0 44252 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_66_475
timestamp 1644511149
transform 1 0 44804 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_66_477
timestamp 1644511149
transform 1 0 44988 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_66_489
timestamp 1644511149
transform 1 0 46092 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_66_512
timestamp 1644511149
transform 1 0 48208 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_3
timestamp 1644511149
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_9
timestamp 1644511149
transform 1 0 1932 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_31
timestamp 1644511149
transform 1 0 3956 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_43
timestamp 1644511149
transform 1 0 5060 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_67_55
timestamp 1644511149
transform 1 0 6164 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_57
timestamp 1644511149
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_69
timestamp 1644511149
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_81
timestamp 1644511149
transform 1 0 8556 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_93
timestamp 1644511149
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_105
timestamp 1644511149
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_111
timestamp 1644511149
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_113
timestamp 1644511149
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_125
timestamp 1644511149
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_137
timestamp 1644511149
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_149
timestamp 1644511149
transform 1 0 14812 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_161
timestamp 1644511149
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_167
timestamp 1644511149
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_169
timestamp 1644511149
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_67_185
timestamp 1644511149
transform 1 0 18124 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_67_193
timestamp 1644511149
transform 1 0 18860 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_67_205
timestamp 1644511149
transform 1 0 19964 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_217
timestamp 1644511149
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_223
timestamp 1644511149
transform 1 0 21620 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_67_225
timestamp 1644511149
transform 1 0 21804 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_233
timestamp 1644511149
transform 1 0 22540 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_67_239
timestamp 1644511149
transform 1 0 23092 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_247
timestamp 1644511149
transform 1 0 23828 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_67_254
timestamp 1644511149
transform 1 0 24472 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_263
timestamp 1644511149
transform 1 0 25300 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_275
timestamp 1644511149
transform 1 0 26404 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_67_279
timestamp 1644511149
transform 1 0 26772 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_67_281
timestamp 1644511149
transform 1 0 26956 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_67_294
timestamp 1644511149
transform 1 0 28152 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_67_314
timestamp 1644511149
transform 1 0 29992 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_67_326
timestamp 1644511149
transform 1 0 31096 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_67_334
timestamp 1644511149
transform 1 0 31832 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_67_337
timestamp 1644511149
transform 1 0 32108 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_349
timestamp 1644511149
transform 1 0 33212 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_361
timestamp 1644511149
transform 1 0 34316 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_373
timestamp 1644511149
transform 1 0 35420 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_385
timestamp 1644511149
transform 1 0 36524 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_391
timestamp 1644511149
transform 1 0 37076 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_393
timestamp 1644511149
transform 1 0 37260 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_405
timestamp 1644511149
transform 1 0 38364 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_417
timestamp 1644511149
transform 1 0 39468 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_429
timestamp 1644511149
transform 1 0 40572 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_67_441
timestamp 1644511149
transform 1 0 41676 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_67_447
timestamp 1644511149
transform 1 0 42228 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_67_449
timestamp 1644511149
transform 1 0 42412 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_461
timestamp 1644511149
transform 1 0 43516 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_473
timestamp 1644511149
transform 1 0 44620 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_67_485
timestamp 1644511149
transform 1 0 45724 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_67_500
timestamp 1644511149
transform 1 0 47104 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_67_505
timestamp 1644511149
transform 1 0 47564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_67_512
timestamp 1644511149
transform 1 0 48208 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_3
timestamp 1644511149
transform 1 0 1380 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_15
timestamp 1644511149
transform 1 0 2484 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_27
timestamp 1644511149
transform 1 0 3588 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_29
timestamp 1644511149
transform 1 0 3772 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_41
timestamp 1644511149
transform 1 0 4876 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_53
timestamp 1644511149
transform 1 0 5980 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_65
timestamp 1644511149
transform 1 0 7084 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_77
timestamp 1644511149
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_83
timestamp 1644511149
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_85
timestamp 1644511149
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_97
timestamp 1644511149
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_109
timestamp 1644511149
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_121
timestamp 1644511149
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_133
timestamp 1644511149
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_139
timestamp 1644511149
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_141
timestamp 1644511149
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_153
timestamp 1644511149
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_68_165
timestamp 1644511149
transform 1 0 16284 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_173
timestamp 1644511149
transform 1 0 17020 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_68_192
timestamp 1644511149
transform 1 0 18768 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_68_205
timestamp 1644511149
transform 1 0 19964 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_68_221
timestamp 1644511149
transform 1 0 21436 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_68_233
timestamp 1644511149
transform 1 0 22540 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_68_242
timestamp 1644511149
transform 1 0 23368 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_68_250
timestamp 1644511149
transform 1 0 24104 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_68_262
timestamp 1644511149
transform 1 0 25208 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_68_270
timestamp 1644511149
transform 1 0 25944 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_68_289
timestamp 1644511149
transform 1 0 27692 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_295
timestamp 1644511149
transform 1 0 28244 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_68_304
timestamp 1644511149
transform 1 0 29072 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_68_313
timestamp 1644511149
transform 1 0 29900 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_325
timestamp 1644511149
transform 1 0 31004 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_337
timestamp 1644511149
transform 1 0 32108 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_349
timestamp 1644511149
transform 1 0 33212 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_68_361
timestamp 1644511149
transform 1 0 34316 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_68_365
timestamp 1644511149
transform 1 0 34684 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_377
timestamp 1644511149
transform 1 0 35788 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_389
timestamp 1644511149
transform 1 0 36892 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_401
timestamp 1644511149
transform 1 0 37996 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_413
timestamp 1644511149
transform 1 0 39100 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_419
timestamp 1644511149
transform 1 0 39652 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_421
timestamp 1644511149
transform 1 0 39836 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_433
timestamp 1644511149
transform 1 0 40940 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_445
timestamp 1644511149
transform 1 0 42044 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_68_457
timestamp 1644511149
transform 1 0 43148 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_68_469
timestamp 1644511149
transform 1 0 44252 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_68_475
timestamp 1644511149
transform 1 0 44804 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_68_477
timestamp 1644511149
transform 1 0 44988 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_68_489
timestamp 1644511149
transform 1 0 46092 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_68_512
timestamp 1644511149
transform 1 0 48208 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_3
timestamp 1644511149
transform 1 0 1380 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_15
timestamp 1644511149
transform 1 0 2484 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_27
timestamp 1644511149
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_39
timestamp 1644511149
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_51
timestamp 1644511149
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_69_55
timestamp 1644511149
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_57
timestamp 1644511149
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_69
timestamp 1644511149
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_81
timestamp 1644511149
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_93
timestamp 1644511149
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_105
timestamp 1644511149
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_111
timestamp 1644511149
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_113
timestamp 1644511149
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_125
timestamp 1644511149
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_137
timestamp 1644511149
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_149
timestamp 1644511149
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_161
timestamp 1644511149
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_167
timestamp 1644511149
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_169
timestamp 1644511149
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_181
timestamp 1644511149
transform 1 0 17756 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_69_191
timestamp 1644511149
transform 1 0 18676 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_211
timestamp 1644511149
transform 1 0 20516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_223
timestamp 1644511149
transform 1 0 21620 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_69_225
timestamp 1644511149
transform 1 0 21804 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_69_233
timestamp 1644511149
transform 1 0 22540 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_69_251
timestamp 1644511149
transform 1 0 24196 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_69_263
timestamp 1644511149
transform 1 0 25300 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_69_273
timestamp 1644511149
transform 1 0 26220 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_279
timestamp 1644511149
transform 1 0 26772 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_69_290
timestamp 1644511149
transform 1 0 27784 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_69_299
timestamp 1644511149
transform 1 0 28612 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_311
timestamp 1644511149
transform 1 0 29716 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_323
timestamp 1644511149
transform 1 0 30820 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_69_335
timestamp 1644511149
transform 1 0 31924 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_337
timestamp 1644511149
transform 1 0 32108 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_349
timestamp 1644511149
transform 1 0 33212 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_361
timestamp 1644511149
transform 1 0 34316 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_373
timestamp 1644511149
transform 1 0 35420 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_385
timestamp 1644511149
transform 1 0 36524 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_391
timestamp 1644511149
transform 1 0 37076 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_393
timestamp 1644511149
transform 1 0 37260 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_405
timestamp 1644511149
transform 1 0 38364 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_417
timestamp 1644511149
transform 1 0 39468 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_429
timestamp 1644511149
transform 1 0 40572 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_69_441
timestamp 1644511149
transform 1 0 41676 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_69_447
timestamp 1644511149
transform 1 0 42228 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_69_449
timestamp 1644511149
transform 1 0 42412 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_461
timestamp 1644511149
transform 1 0 43516 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_473
timestamp 1644511149
transform 1 0 44620 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_69_485
timestamp 1644511149
transform 1 0 45724 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_69_500
timestamp 1644511149
transform 1 0 47104 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_69_508
timestamp 1644511149
transform 1 0 47840 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_70_7
timestamp 1644511149
transform 1 0 1748 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_70_19
timestamp 1644511149
transform 1 0 2852 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_70_27
timestamp 1644511149
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_29
timestamp 1644511149
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_41
timestamp 1644511149
transform 1 0 4876 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_53
timestamp 1644511149
transform 1 0 5980 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_65
timestamp 1644511149
transform 1 0 7084 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_77
timestamp 1644511149
transform 1 0 8188 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_83
timestamp 1644511149
transform 1 0 8740 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_85
timestamp 1644511149
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_97
timestamp 1644511149
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_109
timestamp 1644511149
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_121
timestamp 1644511149
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_133
timestamp 1644511149
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_139
timestamp 1644511149
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_141
timestamp 1644511149
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_153
timestamp 1644511149
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_165
timestamp 1644511149
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_177
timestamp 1644511149
transform 1 0 17388 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_189
timestamp 1644511149
transform 1 0 18492 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_195
timestamp 1644511149
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_70_197
timestamp 1644511149
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_205
timestamp 1644511149
transform 1 0 19964 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_217
timestamp 1644511149
transform 1 0 21068 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_70_229
timestamp 1644511149
transform 1 0 22172 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_70_239
timestamp 1644511149
transform 1 0 23092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_251
timestamp 1644511149
transform 1 0 24196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_70_253
timestamp 1644511149
transform 1 0 24380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_270
timestamp 1644511149
transform 1 0 25944 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_282
timestamp 1644511149
transform 1 0 27048 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_294
timestamp 1644511149
transform 1 0 28152 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_70_306
timestamp 1644511149
transform 1 0 29256 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_70_309
timestamp 1644511149
transform 1 0 29532 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_321
timestamp 1644511149
transform 1 0 30636 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_333
timestamp 1644511149
transform 1 0 31740 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_345
timestamp 1644511149
transform 1 0 32844 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_357
timestamp 1644511149
transform 1 0 33948 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_363
timestamp 1644511149
transform 1 0 34500 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_365
timestamp 1644511149
transform 1 0 34684 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_377
timestamp 1644511149
transform 1 0 35788 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_389
timestamp 1644511149
transform 1 0 36892 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_401
timestamp 1644511149
transform 1 0 37996 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_413
timestamp 1644511149
transform 1 0 39100 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_419
timestamp 1644511149
transform 1 0 39652 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_421
timestamp 1644511149
transform 1 0 39836 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_433
timestamp 1644511149
transform 1 0 40940 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_445
timestamp 1644511149
transform 1 0 42044 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_457
timestamp 1644511149
transform 1 0 43148 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_70_469
timestamp 1644511149
transform 1 0 44252 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_70_475
timestamp 1644511149
transform 1 0 44804 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_70_477
timestamp 1644511149
transform 1 0 44988 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_70_489
timestamp 1644511149
transform 1 0 46092 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_70_501
timestamp 1644511149
transform 1 0 47196 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_70_512
timestamp 1644511149
transform 1 0 48208 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_3
timestamp 1644511149
transform 1 0 1380 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_71_11
timestamp 1644511149
transform 1 0 2116 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_18
timestamp 1644511149
transform 1 0 2760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_30
timestamp 1644511149
transform 1 0 3864 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_42
timestamp 1644511149
transform 1 0 4968 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_71_54
timestamp 1644511149
transform 1 0 6072 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_71_57
timestamp 1644511149
transform 1 0 6348 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_69
timestamp 1644511149
transform 1 0 7452 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_81
timestamp 1644511149
transform 1 0 8556 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_93
timestamp 1644511149
transform 1 0 9660 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_105
timestamp 1644511149
transform 1 0 10764 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_111
timestamp 1644511149
transform 1 0 11316 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_113
timestamp 1644511149
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_125
timestamp 1644511149
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_137
timestamp 1644511149
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_149
timestamp 1644511149
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_161
timestamp 1644511149
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_167
timestamp 1644511149
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_169
timestamp 1644511149
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_181
timestamp 1644511149
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_71_201
timestamp 1644511149
transform 1 0 19596 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_71_211
timestamp 1644511149
transform 1 0 20516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_71_223
timestamp 1644511149
transform 1 0 21620 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_71_233
timestamp 1644511149
transform 1 0 22540 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_239
timestamp 1644511149
transform 1 0 23092 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_256
timestamp 1644511149
transform 1 0 24656 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_268
timestamp 1644511149
transform 1 0 25760 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_281
timestamp 1644511149
transform 1 0 26956 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_293
timestamp 1644511149
transform 1 0 28060 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_305
timestamp 1644511149
transform 1 0 29164 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_317
timestamp 1644511149
transform 1 0 30268 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_329
timestamp 1644511149
transform 1 0 31372 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_335
timestamp 1644511149
transform 1 0 31924 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_337
timestamp 1644511149
transform 1 0 32108 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_349
timestamp 1644511149
transform 1 0 33212 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_361
timestamp 1644511149
transform 1 0 34316 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_373
timestamp 1644511149
transform 1 0 35420 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_385
timestamp 1644511149
transform 1 0 36524 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_391
timestamp 1644511149
transform 1 0 37076 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_393
timestamp 1644511149
transform 1 0 37260 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_405
timestamp 1644511149
transform 1 0 38364 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_417
timestamp 1644511149
transform 1 0 39468 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_429
timestamp 1644511149
transform 1 0 40572 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_71_441
timestamp 1644511149
transform 1 0 41676 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_71_447
timestamp 1644511149
transform 1 0 42228 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_71_449
timestamp 1644511149
transform 1 0 42412 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_461
timestamp 1644511149
transform 1 0 43516 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_71_473
timestamp 1644511149
transform 1 0 44620 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_71_485
timestamp 1644511149
transform 1 0 45724 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_71_493
timestamp 1644511149
transform 1 0 46460 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_71_498
timestamp 1644511149
transform 1 0 46920 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_71_508
timestamp 1644511149
transform 1 0 47840 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_72_24
timestamp 1644511149
transform 1 0 3312 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_72_29
timestamp 1644511149
transform 1 0 3772 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_41
timestamp 1644511149
transform 1 0 4876 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_53
timestamp 1644511149
transform 1 0 5980 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_65
timestamp 1644511149
transform 1 0 7084 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_77
timestamp 1644511149
transform 1 0 8188 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_83
timestamp 1644511149
transform 1 0 8740 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_85
timestamp 1644511149
transform 1 0 8924 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_97
timestamp 1644511149
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_109
timestamp 1644511149
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_121
timestamp 1644511149
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_133
timestamp 1644511149
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_139
timestamp 1644511149
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_141
timestamp 1644511149
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_153
timestamp 1644511149
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_165
timestamp 1644511149
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_177
timestamp 1644511149
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_189
timestamp 1644511149
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_195
timestamp 1644511149
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_72_213
timestamp 1644511149
transform 1 0 20700 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_72_235
timestamp 1644511149
transform 1 0 22724 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_72_247
timestamp 1644511149
transform 1 0 23828 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_72_251
timestamp 1644511149
transform 1 0 24196 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_253
timestamp 1644511149
transform 1 0 24380 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_265
timestamp 1644511149
transform 1 0 25484 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_277
timestamp 1644511149
transform 1 0 26588 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_289
timestamp 1644511149
transform 1 0 27692 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_301
timestamp 1644511149
transform 1 0 28796 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_307
timestamp 1644511149
transform 1 0 29348 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_309
timestamp 1644511149
transform 1 0 29532 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_321
timestamp 1644511149
transform 1 0 30636 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_333
timestamp 1644511149
transform 1 0 31740 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_345
timestamp 1644511149
transform 1 0 32844 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_357
timestamp 1644511149
transform 1 0 33948 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_363
timestamp 1644511149
transform 1 0 34500 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_365
timestamp 1644511149
transform 1 0 34684 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_377
timestamp 1644511149
transform 1 0 35788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_389
timestamp 1644511149
transform 1 0 36892 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_401
timestamp 1644511149
transform 1 0 37996 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_413
timestamp 1644511149
transform 1 0 39100 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_419
timestamp 1644511149
transform 1 0 39652 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_421
timestamp 1644511149
transform 1 0 39836 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_433
timestamp 1644511149
transform 1 0 40940 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_445
timestamp 1644511149
transform 1 0 42044 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_72_457
timestamp 1644511149
transform 1 0 43148 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_72_469
timestamp 1644511149
transform 1 0 44252 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_72_475
timestamp 1644511149
transform 1 0 44804 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_72_477
timestamp 1644511149
transform 1 0 44988 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_72_489
timestamp 1644511149
transform 1 0 46092 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_72_512
timestamp 1644511149
transform 1 0 48208 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_73_3
timestamp 1644511149
transform 1 0 1380 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_7
timestamp 1644511149
transform 1 0 1748 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_11
timestamp 1644511149
transform 1 0 2116 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_23
timestamp 1644511149
transform 1 0 3220 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_35
timestamp 1644511149
transform 1 0 4324 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_73_47
timestamp 1644511149
transform 1 0 5428 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_73_55
timestamp 1644511149
transform 1 0 6164 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_57
timestamp 1644511149
transform 1 0 6348 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_69
timestamp 1644511149
transform 1 0 7452 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_81
timestamp 1644511149
transform 1 0 8556 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_93
timestamp 1644511149
transform 1 0 9660 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_105
timestamp 1644511149
transform 1 0 10764 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_111
timestamp 1644511149
transform 1 0 11316 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_113
timestamp 1644511149
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_125
timestamp 1644511149
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_137
timestamp 1644511149
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_149
timestamp 1644511149
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_161
timestamp 1644511149
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_167
timestamp 1644511149
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_169
timestamp 1644511149
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_181
timestamp 1644511149
transform 1 0 17756 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_193
timestamp 1644511149
transform 1 0 18860 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_205
timestamp 1644511149
transform 1 0 19964 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_217
timestamp 1644511149
transform 1 0 21068 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_223
timestamp 1644511149
transform 1 0 21620 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_73_225
timestamp 1644511149
transform 1 0 21804 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_73_239
timestamp 1644511149
transform 1 0 23092 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_251
timestamp 1644511149
transform 1 0 24196 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_263
timestamp 1644511149
transform 1 0 25300 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_73_275
timestamp 1644511149
transform 1 0 26404 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_73_279
timestamp 1644511149
transform 1 0 26772 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_281
timestamp 1644511149
transform 1 0 26956 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_293
timestamp 1644511149
transform 1 0 28060 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_305
timestamp 1644511149
transform 1 0 29164 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_317
timestamp 1644511149
transform 1 0 30268 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_329
timestamp 1644511149
transform 1 0 31372 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_335
timestamp 1644511149
transform 1 0 31924 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_337
timestamp 1644511149
transform 1 0 32108 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_349
timestamp 1644511149
transform 1 0 33212 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_361
timestamp 1644511149
transform 1 0 34316 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_373
timestamp 1644511149
transform 1 0 35420 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_385
timestamp 1644511149
transform 1 0 36524 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_391
timestamp 1644511149
transform 1 0 37076 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_393
timestamp 1644511149
transform 1 0 37260 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_405
timestamp 1644511149
transform 1 0 38364 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_417
timestamp 1644511149
transform 1 0 39468 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_429
timestamp 1644511149
transform 1 0 40572 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_441
timestamp 1644511149
transform 1 0 41676 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_447
timestamp 1644511149
transform 1 0 42228 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_73_449
timestamp 1644511149
transform 1 0 42412 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_461
timestamp 1644511149
transform 1 0 43516 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_473
timestamp 1644511149
transform 1 0 44620 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_73_485
timestamp 1644511149
transform 1 0 45724 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_73_497
timestamp 1644511149
transform 1 0 46828 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_73_503
timestamp 1644511149
transform 1 0 47380 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_73_512
timestamp 1644511149
transform 1 0 48208 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_74_3
timestamp 1644511149
transform 1 0 1380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_15
timestamp 1644511149
transform 1 0 2484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_74_27
timestamp 1644511149
transform 1 0 3588 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_29
timestamp 1644511149
transform 1 0 3772 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_41
timestamp 1644511149
transform 1 0 4876 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_53
timestamp 1644511149
transform 1 0 5980 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_65
timestamp 1644511149
transform 1 0 7084 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_77
timestamp 1644511149
transform 1 0 8188 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_83
timestamp 1644511149
transform 1 0 8740 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_85
timestamp 1644511149
transform 1 0 8924 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_97
timestamp 1644511149
transform 1 0 10028 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_109
timestamp 1644511149
transform 1 0 11132 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_121
timestamp 1644511149
transform 1 0 12236 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_133
timestamp 1644511149
transform 1 0 13340 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_139
timestamp 1644511149
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_141
timestamp 1644511149
transform 1 0 14076 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_153
timestamp 1644511149
transform 1 0 15180 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_165
timestamp 1644511149
transform 1 0 16284 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_177
timestamp 1644511149
transform 1 0 17388 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_189
timestamp 1644511149
transform 1 0 18492 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_195
timestamp 1644511149
transform 1 0 19044 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_197
timestamp 1644511149
transform 1 0 19228 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_209
timestamp 1644511149
transform 1 0 20332 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_221
timestamp 1644511149
transform 1 0 21436 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_233
timestamp 1644511149
transform 1 0 22540 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_245
timestamp 1644511149
transform 1 0 23644 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_251
timestamp 1644511149
transform 1 0 24196 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_253
timestamp 1644511149
transform 1 0 24380 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_265
timestamp 1644511149
transform 1 0 25484 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_277
timestamp 1644511149
transform 1 0 26588 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_289
timestamp 1644511149
transform 1 0 27692 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_301
timestamp 1644511149
transform 1 0 28796 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_307
timestamp 1644511149
transform 1 0 29348 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_309
timestamp 1644511149
transform 1 0 29532 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_321
timestamp 1644511149
transform 1 0 30636 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_333
timestamp 1644511149
transform 1 0 31740 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_345
timestamp 1644511149
transform 1 0 32844 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_357
timestamp 1644511149
transform 1 0 33948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_363
timestamp 1644511149
transform 1 0 34500 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_365
timestamp 1644511149
transform 1 0 34684 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_377
timestamp 1644511149
transform 1 0 35788 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_389
timestamp 1644511149
transform 1 0 36892 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_401
timestamp 1644511149
transform 1 0 37996 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_413
timestamp 1644511149
transform 1 0 39100 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_419
timestamp 1644511149
transform 1 0 39652 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_421
timestamp 1644511149
transform 1 0 39836 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_433
timestamp 1644511149
transform 1 0 40940 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_445
timestamp 1644511149
transform 1 0 42044 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_74_457
timestamp 1644511149
transform 1 0 43148 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_74_469
timestamp 1644511149
transform 1 0 44252 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_74_475
timestamp 1644511149
transform 1 0 44804 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_74_477
timestamp 1644511149
transform 1 0 44988 0 1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_74_489
timestamp 1644511149
transform 1 0 46092 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_74_512
timestamp 1644511149
transform 1 0 48208 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_75_3
timestamp 1644511149
transform 1 0 1380 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_15
timestamp 1644511149
transform 1 0 2484 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_27
timestamp 1644511149
transform 1 0 3588 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_39
timestamp 1644511149
transform 1 0 4692 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_51
timestamp 1644511149
transform 1 0 5796 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_75_55
timestamp 1644511149
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_57
timestamp 1644511149
transform 1 0 6348 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_69
timestamp 1644511149
transform 1 0 7452 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_81
timestamp 1644511149
transform 1 0 8556 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_93
timestamp 1644511149
transform 1 0 9660 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_105
timestamp 1644511149
transform 1 0 10764 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_111
timestamp 1644511149
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_113
timestamp 1644511149
transform 1 0 11500 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_125
timestamp 1644511149
transform 1 0 12604 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_137
timestamp 1644511149
transform 1 0 13708 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_149
timestamp 1644511149
transform 1 0 14812 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_161
timestamp 1644511149
transform 1 0 15916 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_167
timestamp 1644511149
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_169
timestamp 1644511149
transform 1 0 16652 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_181
timestamp 1644511149
transform 1 0 17756 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_193
timestamp 1644511149
transform 1 0 18860 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_205
timestamp 1644511149
transform 1 0 19964 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_217
timestamp 1644511149
transform 1 0 21068 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_223
timestamp 1644511149
transform 1 0 21620 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_225
timestamp 1644511149
transform 1 0 21804 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_237
timestamp 1644511149
transform 1 0 22908 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_249
timestamp 1644511149
transform 1 0 24012 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_261
timestamp 1644511149
transform 1 0 25116 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_273
timestamp 1644511149
transform 1 0 26220 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_279
timestamp 1644511149
transform 1 0 26772 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_281
timestamp 1644511149
transform 1 0 26956 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_293
timestamp 1644511149
transform 1 0 28060 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_305
timestamp 1644511149
transform 1 0 29164 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_317
timestamp 1644511149
transform 1 0 30268 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_329
timestamp 1644511149
transform 1 0 31372 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_335
timestamp 1644511149
transform 1 0 31924 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_337
timestamp 1644511149
transform 1 0 32108 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_349
timestamp 1644511149
transform 1 0 33212 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_361
timestamp 1644511149
transform 1 0 34316 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_373
timestamp 1644511149
transform 1 0 35420 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_385
timestamp 1644511149
transform 1 0 36524 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_391
timestamp 1644511149
transform 1 0 37076 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_393
timestamp 1644511149
transform 1 0 37260 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_405
timestamp 1644511149
transform 1 0 38364 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_417
timestamp 1644511149
transform 1 0 39468 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_429
timestamp 1644511149
transform 1 0 40572 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_75_441
timestamp 1644511149
transform 1 0 41676 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_75_447
timestamp 1644511149
transform 1 0 42228 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_75_449
timestamp 1644511149
transform 1 0 42412 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_461
timestamp 1644511149
transform 1 0 43516 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_473
timestamp 1644511149
transform 1 0 44620 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_75_485
timestamp 1644511149
transform 1 0 45724 0 -1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_75_500
timestamp 1644511149
transform 1 0 47104 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_75_505
timestamp 1644511149
transform 1 0 47564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_75_512
timestamp 1644511149
transform 1 0 48208 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_3
timestamp 1644511149
transform 1 0 1380 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_13
timestamp 1644511149
transform 1 0 2300 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_76_20
timestamp 1644511149
transform 1 0 2944 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_29
timestamp 1644511149
transform 1 0 3772 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_41
timestamp 1644511149
transform 1 0 4876 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_53
timestamp 1644511149
transform 1 0 5980 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_65
timestamp 1644511149
transform 1 0 7084 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_77
timestamp 1644511149
transform 1 0 8188 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_83
timestamp 1644511149
transform 1 0 8740 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_85
timestamp 1644511149
transform 1 0 8924 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_97
timestamp 1644511149
transform 1 0 10028 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_109
timestamp 1644511149
transform 1 0 11132 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_121
timestamp 1644511149
transform 1 0 12236 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_133
timestamp 1644511149
transform 1 0 13340 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_139
timestamp 1644511149
transform 1 0 13892 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_141
timestamp 1644511149
transform 1 0 14076 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_153
timestamp 1644511149
transform 1 0 15180 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_165
timestamp 1644511149
transform 1 0 16284 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_177
timestamp 1644511149
transform 1 0 17388 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_189
timestamp 1644511149
transform 1 0 18492 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_195
timestamp 1644511149
transform 1 0 19044 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_197
timestamp 1644511149
transform 1 0 19228 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_209
timestamp 1644511149
transform 1 0 20332 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_221
timestamp 1644511149
transform 1 0 21436 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_233
timestamp 1644511149
transform 1 0 22540 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_245
timestamp 1644511149
transform 1 0 23644 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_251
timestamp 1644511149
transform 1 0 24196 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_253
timestamp 1644511149
transform 1 0 24380 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_265
timestamp 1644511149
transform 1 0 25484 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_277
timestamp 1644511149
transform 1 0 26588 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_283
timestamp 1644511149
transform 1 0 27140 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_76_300
timestamp 1644511149
transform 1 0 28704 0 1 43520
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_76_309
timestamp 1644511149
transform 1 0 29532 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_321
timestamp 1644511149
transform 1 0 30636 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_333
timestamp 1644511149
transform 1 0 31740 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_345
timestamp 1644511149
transform 1 0 32844 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_357
timestamp 1644511149
transform 1 0 33948 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_363
timestamp 1644511149
transform 1 0 34500 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_365
timestamp 1644511149
transform 1 0 34684 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_377
timestamp 1644511149
transform 1 0 35788 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_389
timestamp 1644511149
transform 1 0 36892 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_401
timestamp 1644511149
transform 1 0 37996 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_413
timestamp 1644511149
transform 1 0 39100 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_419
timestamp 1644511149
transform 1 0 39652 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_421
timestamp 1644511149
transform 1 0 39836 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_433
timestamp 1644511149
transform 1 0 40940 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_445
timestamp 1644511149
transform 1 0 42044 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_76_457
timestamp 1644511149
transform 1 0 43148 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_76_469
timestamp 1644511149
transform 1 0 44252 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_76_475
timestamp 1644511149
transform 1 0 44804 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_76_477
timestamp 1644511149
transform 1 0 44988 0 1 43520
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_76_489
timestamp 1644511149
transform 1 0 46092 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_76_493
timestamp 1644511149
transform 1 0 46460 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_76_497
timestamp 1644511149
transform 1 0 46828 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_504
timestamp 1644511149
transform 1 0 47472 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_76_512
timestamp 1644511149
transform 1 0 48208 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_3
timestamp 1644511149
transform 1 0 1380 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_13
timestamp 1644511149
transform 1 0 2300 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_20
timestamp 1644511149
transform 1 0 2944 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_77_27
timestamp 1644511149
transform 1 0 3588 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_39
timestamp 1644511149
transform 1 0 4692 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_51
timestamp 1644511149
transform 1 0 5796 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_55
timestamp 1644511149
transform 1 0 6164 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_57
timestamp 1644511149
transform 1 0 6348 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_69
timestamp 1644511149
transform 1 0 7452 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_81
timestamp 1644511149
transform 1 0 8556 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_93
timestamp 1644511149
transform 1 0 9660 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_105
timestamp 1644511149
transform 1 0 10764 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_111
timestamp 1644511149
transform 1 0 11316 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_113
timestamp 1644511149
transform 1 0 11500 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_125
timestamp 1644511149
transform 1 0 12604 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_137
timestamp 1644511149
transform 1 0 13708 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_149
timestamp 1644511149
transform 1 0 14812 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_161
timestamp 1644511149
transform 1 0 15916 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_167
timestamp 1644511149
transform 1 0 16468 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_169
timestamp 1644511149
transform 1 0 16652 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_181
timestamp 1644511149
transform 1 0 17756 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_193
timestamp 1644511149
transform 1 0 18860 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_205
timestamp 1644511149
transform 1 0 19964 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_217
timestamp 1644511149
transform 1 0 21068 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_223
timestamp 1644511149
transform 1 0 21620 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_225
timestamp 1644511149
transform 1 0 21804 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_237
timestamp 1644511149
transform 1 0 22908 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_249
timestamp 1644511149
transform 1 0 24012 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_261
timestamp 1644511149
transform 1 0 25116 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_273
timestamp 1644511149
transform 1 0 26220 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_279
timestamp 1644511149
transform 1 0 26772 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_281
timestamp 1644511149
transform 1 0 26956 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_293
timestamp 1644511149
transform 1 0 28060 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_305
timestamp 1644511149
transform 1 0 29164 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_317
timestamp 1644511149
transform 1 0 30268 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_329
timestamp 1644511149
transform 1 0 31372 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_335
timestamp 1644511149
transform 1 0 31924 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_337
timestamp 1644511149
transform 1 0 32108 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_349
timestamp 1644511149
transform 1 0 33212 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_361
timestamp 1644511149
transform 1 0 34316 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_373
timestamp 1644511149
transform 1 0 35420 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_385
timestamp 1644511149
transform 1 0 36524 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_391
timestamp 1644511149
transform 1 0 37076 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_393
timestamp 1644511149
transform 1 0 37260 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_405
timestamp 1644511149
transform 1 0 38364 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_417
timestamp 1644511149
transform 1 0 39468 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_429
timestamp 1644511149
transform 1 0 40572 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_77_441
timestamp 1644511149
transform 1 0 41676 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_77_447
timestamp 1644511149
transform 1 0 42228 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_77_449
timestamp 1644511149
transform 1 0 42412 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_77_461
timestamp 1644511149
transform 1 0 43516 0 -1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_77_473
timestamp 1644511149
transform 1 0 44620 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_77_477
timestamp 1644511149
transform 1 0 44988 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_77_481
timestamp 1644511149
transform 1 0 45356 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_77_489
timestamp 1644511149
transform 1 0 46092 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_77_493
timestamp 1644511149
transform 1 0 46460 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_77_500
timestamp 1644511149
transform 1 0 47104 0 -1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_77_508
timestamp 1644511149
transform 1 0 47840 0 -1 44608
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_78_24
timestamp 1644511149
transform 1 0 3312 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_78_29
timestamp 1644511149
transform 1 0 3772 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_41
timestamp 1644511149
transform 1 0 4876 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_53
timestamp 1644511149
transform 1 0 5980 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_65
timestamp 1644511149
transform 1 0 7084 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_77
timestamp 1644511149
transform 1 0 8188 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_83
timestamp 1644511149
transform 1 0 8740 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_85
timestamp 1644511149
transform 1 0 8924 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_97
timestamp 1644511149
transform 1 0 10028 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_109
timestamp 1644511149
transform 1 0 11132 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_121
timestamp 1644511149
transform 1 0 12236 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_133
timestamp 1644511149
transform 1 0 13340 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_139
timestamp 1644511149
transform 1 0 13892 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_141
timestamp 1644511149
transform 1 0 14076 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_153
timestamp 1644511149
transform 1 0 15180 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_165
timestamp 1644511149
transform 1 0 16284 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_177
timestamp 1644511149
transform 1 0 17388 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_189
timestamp 1644511149
transform 1 0 18492 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_195
timestamp 1644511149
transform 1 0 19044 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_197
timestamp 1644511149
transform 1 0 19228 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_209
timestamp 1644511149
transform 1 0 20332 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_221
timestamp 1644511149
transform 1 0 21436 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_233
timestamp 1644511149
transform 1 0 22540 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_245
timestamp 1644511149
transform 1 0 23644 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_251
timestamp 1644511149
transform 1 0 24196 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_253
timestamp 1644511149
transform 1 0 24380 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_265
timestamp 1644511149
transform 1 0 25484 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_277
timestamp 1644511149
transform 1 0 26588 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_289
timestamp 1644511149
transform 1 0 27692 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_301
timestamp 1644511149
transform 1 0 28796 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_307
timestamp 1644511149
transform 1 0 29348 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_309
timestamp 1644511149
transform 1 0 29532 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_321
timestamp 1644511149
transform 1 0 30636 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_333
timestamp 1644511149
transform 1 0 31740 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_345
timestamp 1644511149
transform 1 0 32844 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_357
timestamp 1644511149
transform 1 0 33948 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_363
timestamp 1644511149
transform 1 0 34500 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_365
timestamp 1644511149
transform 1 0 34684 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_377
timestamp 1644511149
transform 1 0 35788 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_389
timestamp 1644511149
transform 1 0 36892 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_401
timestamp 1644511149
transform 1 0 37996 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_413
timestamp 1644511149
transform 1 0 39100 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_419
timestamp 1644511149
transform 1 0 39652 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_78_421
timestamp 1644511149
transform 1 0 39836 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_433
timestamp 1644511149
transform 1 0 40940 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_445
timestamp 1644511149
transform 1 0 42044 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_78_457
timestamp 1644511149
transform 1 0 43148 0 1 44608
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_78_469
timestamp 1644511149
transform 1 0 44252 0 1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_78_475
timestamp 1644511149
transform 1 0 44804 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_78_480
timestamp 1644511149
transform 1 0 45264 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_487
timestamp 1644511149
transform 1 0 45908 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_78_512
timestamp 1644511149
transform 1 0 48208 0 1 44608
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_3
timestamp 1644511149
transform 1 0 1380 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_28
timestamp 1644511149
transform 1 0 3680 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_40
timestamp 1644511149
transform 1 0 4784 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_52
timestamp 1644511149
transform 1 0 5888 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_79_57
timestamp 1644511149
transform 1 0 6348 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_69
timestamp 1644511149
transform 1 0 7452 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_81
timestamp 1644511149
transform 1 0 8556 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_93
timestamp 1644511149
transform 1 0 9660 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_105
timestamp 1644511149
transform 1 0 10764 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_111
timestamp 1644511149
transform 1 0 11316 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_113
timestamp 1644511149
transform 1 0 11500 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_125
timestamp 1644511149
transform 1 0 12604 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_137
timestamp 1644511149
transform 1 0 13708 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_149
timestamp 1644511149
transform 1 0 14812 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_161
timestamp 1644511149
transform 1 0 15916 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_167
timestamp 1644511149
transform 1 0 16468 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_169
timestamp 1644511149
transform 1 0 16652 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_181
timestamp 1644511149
transform 1 0 17756 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_193
timestamp 1644511149
transform 1 0 18860 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_205
timestamp 1644511149
transform 1 0 19964 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_217
timestamp 1644511149
transform 1 0 21068 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_223
timestamp 1644511149
transform 1 0 21620 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_225
timestamp 1644511149
transform 1 0 21804 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_237
timestamp 1644511149
transform 1 0 22908 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_249
timestamp 1644511149
transform 1 0 24012 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_261
timestamp 1644511149
transform 1 0 25116 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_273
timestamp 1644511149
transform 1 0 26220 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_279
timestamp 1644511149
transform 1 0 26772 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_281
timestamp 1644511149
transform 1 0 26956 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_293
timestamp 1644511149
transform 1 0 28060 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_305
timestamp 1644511149
transform 1 0 29164 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_317
timestamp 1644511149
transform 1 0 30268 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_329
timestamp 1644511149
transform 1 0 31372 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_335
timestamp 1644511149
transform 1 0 31924 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_337
timestamp 1644511149
transform 1 0 32108 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_349
timestamp 1644511149
transform 1 0 33212 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_361
timestamp 1644511149
transform 1 0 34316 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_373
timestamp 1644511149
transform 1 0 35420 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_385
timestamp 1644511149
transform 1 0 36524 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_391
timestamp 1644511149
transform 1 0 37076 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_393
timestamp 1644511149
transform 1 0 37260 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_405
timestamp 1644511149
transform 1 0 38364 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_417
timestamp 1644511149
transform 1 0 39468 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_79_429
timestamp 1644511149
transform 1 0 40572 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_79_441
timestamp 1644511149
transform 1 0 41676 0 -1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_79_447
timestamp 1644511149
transform 1 0 42228 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_79_449
timestamp 1644511149
transform 1 0 42412 0 -1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_79_461
timestamp 1644511149
transform 1 0 43516 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_468
timestamp 1644511149
transform 1 0 44160 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_475
timestamp 1644511149
transform 1 0 44804 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_79_500
timestamp 1644511149
transform 1 0 47104 0 -1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_79_508
timestamp 1644511149
transform 1 0 47840 0 -1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_80_7
timestamp 1644511149
transform 1 0 1748 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_80_16
timestamp 1644511149
transform 1 0 2576 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_23
timestamp 1644511149
transform 1 0 3220 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_80_27
timestamp 1644511149
transform 1 0 3588 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_32
timestamp 1644511149
transform 1 0 4048 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_44
timestamp 1644511149
transform 1 0 5152 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_56
timestamp 1644511149
transform 1 0 6256 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_68
timestamp 1644511149
transform 1 0 7360 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_80_80
timestamp 1644511149
transform 1 0 8464 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_80_85
timestamp 1644511149
transform 1 0 8924 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_97
timestamp 1644511149
transform 1 0 10028 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_109
timestamp 1644511149
transform 1 0 11132 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_121
timestamp 1644511149
transform 1 0 12236 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_133
timestamp 1644511149
transform 1 0 13340 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_139
timestamp 1644511149
transform 1 0 13892 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_141
timestamp 1644511149
transform 1 0 14076 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_153
timestamp 1644511149
transform 1 0 15180 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_165
timestamp 1644511149
transform 1 0 16284 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_177
timestamp 1644511149
transform 1 0 17388 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_189
timestamp 1644511149
transform 1 0 18492 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_195
timestamp 1644511149
transform 1 0 19044 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_197
timestamp 1644511149
transform 1 0 19228 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_209
timestamp 1644511149
transform 1 0 20332 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_221
timestamp 1644511149
transform 1 0 21436 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_233
timestamp 1644511149
transform 1 0 22540 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_245
timestamp 1644511149
transform 1 0 23644 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_251
timestamp 1644511149
transform 1 0 24196 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_253
timestamp 1644511149
transform 1 0 24380 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_265
timestamp 1644511149
transform 1 0 25484 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_277
timestamp 1644511149
transform 1 0 26588 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_289
timestamp 1644511149
transform 1 0 27692 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_301
timestamp 1644511149
transform 1 0 28796 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_307
timestamp 1644511149
transform 1 0 29348 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_309
timestamp 1644511149
transform 1 0 29532 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_321
timestamp 1644511149
transform 1 0 30636 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_333
timestamp 1644511149
transform 1 0 31740 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_345
timestamp 1644511149
transform 1 0 32844 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_357
timestamp 1644511149
transform 1 0 33948 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_363
timestamp 1644511149
transform 1 0 34500 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_365
timestamp 1644511149
transform 1 0 34684 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_377
timestamp 1644511149
transform 1 0 35788 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_389
timestamp 1644511149
transform 1 0 36892 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_80_401
timestamp 1644511149
transform 1 0 37996 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_80_413
timestamp 1644511149
transform 1 0 39100 0 1 45696
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_80_419
timestamp 1644511149
transform 1 0 39652 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_80_421
timestamp 1644511149
transform 1 0 39836 0 1 45696
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_80_433
timestamp 1644511149
transform 1 0 40940 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_80_441
timestamp 1644511149
transform 1 0 41676 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_80_445
timestamp 1644511149
transform 1 0 42044 0 1 45696
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_80_451
timestamp 1644511149
transform 1 0 42596 0 1 45696
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_80_459
timestamp 1644511149
transform 1 0 43332 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_80_465
timestamp 1644511149
transform 1 0 43884 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_472
timestamp 1644511149
transform 1 0 44528 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_480
timestamp 1644511149
transform 1 0 45264 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_487
timestamp 1644511149
transform 1 0 45908 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_80_512
timestamp 1644511149
transform 1 0 48208 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_6
timestamp 1644511149
transform 1 0 1656 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_14
timestamp 1644511149
transform 1 0 2392 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_21
timestamp 1644511149
transform 1 0 3036 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_81_28
timestamp 1644511149
transform 1 0 3680 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_81_35
timestamp 1644511149
transform 1 0 4324 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_43
timestamp 1644511149
transform 1 0 5060 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_47
timestamp 1644511149
transform 1 0 5428 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_81_55
timestamp 1644511149
transform 1 0 6164 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_57
timestamp 1644511149
transform 1 0 6348 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_69
timestamp 1644511149
transform 1 0 7452 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_81
timestamp 1644511149
transform 1 0 8556 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_93
timestamp 1644511149
transform 1 0 9660 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_105
timestamp 1644511149
transform 1 0 10764 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_111
timestamp 1644511149
transform 1 0 11316 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_113
timestamp 1644511149
transform 1 0 11500 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_125
timestamp 1644511149
transform 1 0 12604 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_137
timestamp 1644511149
transform 1 0 13708 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_149
timestamp 1644511149
transform 1 0 14812 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_161
timestamp 1644511149
transform 1 0 15916 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_167
timestamp 1644511149
transform 1 0 16468 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_169
timestamp 1644511149
transform 1 0 16652 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_181
timestamp 1644511149
transform 1 0 17756 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_193
timestamp 1644511149
transform 1 0 18860 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_205
timestamp 1644511149
transform 1 0 19964 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_217
timestamp 1644511149
transform 1 0 21068 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_223
timestamp 1644511149
transform 1 0 21620 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_225
timestamp 1644511149
transform 1 0 21804 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_237
timestamp 1644511149
transform 1 0 22908 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_249
timestamp 1644511149
transform 1 0 24012 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_261
timestamp 1644511149
transform 1 0 25116 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_273
timestamp 1644511149
transform 1 0 26220 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_279
timestamp 1644511149
transform 1 0 26772 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_281
timestamp 1644511149
transform 1 0 26956 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_293
timestamp 1644511149
transform 1 0 28060 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_305
timestamp 1644511149
transform 1 0 29164 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_317
timestamp 1644511149
transform 1 0 30268 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_329
timestamp 1644511149
transform 1 0 31372 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_335
timestamp 1644511149
transform 1 0 31924 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_337
timestamp 1644511149
transform 1 0 32108 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_349
timestamp 1644511149
transform 1 0 33212 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_361
timestamp 1644511149
transform 1 0 34316 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_373
timestamp 1644511149
transform 1 0 35420 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_385
timestamp 1644511149
transform 1 0 36524 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_391
timestamp 1644511149
transform 1 0 37076 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_81_393
timestamp 1644511149
transform 1 0 37260 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_405
timestamp 1644511149
transform 1 0 38364 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_417
timestamp 1644511149
transform 1 0 39468 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_81_429
timestamp 1644511149
transform 1 0 40572 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_81_441
timestamp 1644511149
transform 1 0 41676 0 -1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_81_447
timestamp 1644511149
transform 1 0 42228 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_81_461
timestamp 1644511149
transform 1 0 43516 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_81_465
timestamp 1644511149
transform 1 0 43884 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_81_469
timestamp 1644511149
transform 1 0 44252 0 -1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_81_477
timestamp 1644511149
transform 1 0 44988 0 -1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_81_500
timestamp 1644511149
transform 1 0 47104 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_81_505
timestamp 1644511149
transform 1 0 47564 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_81_512
timestamp 1644511149
transform 1 0 48208 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_24
timestamp 1644511149
transform 1 0 3312 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_32
timestamp 1644511149
transform 1 0 4048 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_38
timestamp 1644511149
transform 1 0 4600 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_42
timestamp 1644511149
transform 1 0 4968 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_49
timestamp 1644511149
transform 1 0 5612 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_58
timestamp 1644511149
transform 1 0 6440 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_65
timestamp 1644511149
transform 1 0 7084 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_71
timestamp 1644511149
transform 1 0 7636 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_82_75
timestamp 1644511149
transform 1 0 8004 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_82_83
timestamp 1644511149
transform 1 0 8740 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_85
timestamp 1644511149
transform 1 0 8924 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_97
timestamp 1644511149
transform 1 0 10028 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_109
timestamp 1644511149
transform 1 0 11132 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_121
timestamp 1644511149
transform 1 0 12236 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_133
timestamp 1644511149
transform 1 0 13340 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_139
timestamp 1644511149
transform 1 0 13892 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_141
timestamp 1644511149
transform 1 0 14076 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_153
timestamp 1644511149
transform 1 0 15180 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_165
timestamp 1644511149
transform 1 0 16284 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_177
timestamp 1644511149
transform 1 0 17388 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_189
timestamp 1644511149
transform 1 0 18492 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_195
timestamp 1644511149
transform 1 0 19044 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_197
timestamp 1644511149
transform 1 0 19228 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_230
timestamp 1644511149
transform 1 0 22264 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_82_242
timestamp 1644511149
transform 1 0 23368 0 1 46784
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_82_250
timestamp 1644511149
transform 1 0 24104 0 1 46784
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_82_253
timestamp 1644511149
transform 1 0 24380 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_265
timestamp 1644511149
transform 1 0 25484 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_277
timestamp 1644511149
transform 1 0 26588 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_82_289
timestamp 1644511149
transform 1 0 27692 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_293
timestamp 1644511149
transform 1 0 28060 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_82_305
timestamp 1644511149
transform 1 0 29164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_82_309
timestamp 1644511149
transform 1 0 29532 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_321
timestamp 1644511149
transform 1 0 30636 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_333
timestamp 1644511149
transform 1 0 31740 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_345
timestamp 1644511149
transform 1 0 32844 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_357
timestamp 1644511149
transform 1 0 33948 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_363
timestamp 1644511149
transform 1 0 34500 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_365
timestamp 1644511149
transform 1 0 34684 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_377
timestamp 1644511149
transform 1 0 35788 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_389
timestamp 1644511149
transform 1 0 36892 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_82_401
timestamp 1644511149
transform 1 0 37996 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_82_413
timestamp 1644511149
transform 1 0 39100 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_82_419
timestamp 1644511149
transform 1 0 39652 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_82_421
timestamp 1644511149
transform 1 0 39836 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_82_433
timestamp 1644511149
transform 1 0 40940 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_82_437
timestamp 1644511149
transform 1 0 41308 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_82_454
timestamp 1644511149
transform 1 0 42872 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_82_470
timestamp 1644511149
transform 1 0 44344 0 1 46784
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_82_480
timestamp 1644511149
transform 1 0 45264 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_487
timestamp 1644511149
transform 1 0 45908 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_82_512
timestamp 1644511149
transform 1 0 48208 0 1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_3
timestamp 1644511149
transform 1 0 1380 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_83_30
timestamp 1644511149
transform 1 0 3864 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_37
timestamp 1644511149
transform 1 0 4508 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_44
timestamp 1644511149
transform 1 0 5152 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_52
timestamp 1644511149
transform 1 0 5888 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_78
timestamp 1644511149
transform 1 0 8280 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_85
timestamp 1644511149
transform 1 0 8924 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_93
timestamp 1644511149
transform 1 0 9660 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_97
timestamp 1644511149
transform 1 0 10028 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_104
timestamp 1644511149
transform 1 0 10672 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_83_113
timestamp 1644511149
transform 1 0 11500 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_125
timestamp 1644511149
transform 1 0 12604 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_83_137
timestamp 1644511149
transform 1 0 13708 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_83_146
timestamp 1644511149
transform 1 0 14536 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_83_158
timestamp 1644511149
transform 1 0 15640 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_166
timestamp 1644511149
transform 1 0 16376 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_172
timestamp 1644511149
transform 1 0 16928 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_179
timestamp 1644511149
transform 1 0 17572 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_191
timestamp 1644511149
transform 1 0 18676 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_203
timestamp 1644511149
transform 1 0 19780 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_210
timestamp 1644511149
transform 1 0 20424 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_83_217
timestamp 1644511149
transform 1 0 21068 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_83_223
timestamp 1644511149
transform 1 0 21620 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_225
timestamp 1644511149
transform 1 0 21804 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_232
timestamp 1644511149
transform 1 0 22448 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_244
timestamp 1644511149
transform 1 0 23552 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_256
timestamp 1644511149
transform 1 0 24656 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_268
timestamp 1644511149
transform 1 0 25760 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_272
timestamp 1644511149
transform 1 0 26128 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_276
timestamp 1644511149
transform 1 0 26496 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_281
timestamp 1644511149
transform 1 0 26956 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_288
timestamp 1644511149
transform 1 0 27600 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_313
timestamp 1644511149
transform 1 0 29900 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_320
timestamp 1644511149
transform 1 0 30544 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_324
timestamp 1644511149
transform 1 0 30912 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_83_328
timestamp 1644511149
transform 1 0 31280 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_83_337
timestamp 1644511149
transform 1 0 32108 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_83_343
timestamp 1644511149
transform 1 0 32660 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_83_351
timestamp 1644511149
transform 1 0 33396 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_373
timestamp 1644511149
transform 1 0 35420 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_83_380
timestamp 1644511149
transform 1 0 36064 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_393
timestamp 1644511149
transform 1 0 37260 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_405
timestamp 1644511149
transform 1 0 38364 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_83_417
timestamp 1644511149
transform 1 0 39468 0 -1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_83_429
timestamp 1644511149
transform 1 0 40572 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_433
timestamp 1644511149
transform 1 0 40940 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_437
timestamp 1644511149
transform 1 0 41308 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_444
timestamp 1644511149
transform 1 0 41952 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_83_458
timestamp 1644511149
transform 1 0 43240 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_83_468
timestamp 1644511149
transform 1 0 44160 0 -1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_83_476
timestamp 1644511149
transform 1 0 44896 0 -1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_83_499
timestamp 1644511149
transform 1 0 47012 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_83_503
timestamp 1644511149
transform 1 0 47380 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_83_505
timestamp 1644511149
transform 1 0 47564 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_83_512
timestamp 1644511149
transform 1 0 48208 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_24
timestamp 1644511149
transform 1 0 3312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_33
timestamp 1644511149
transform 1 0 4140 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_58
timestamp 1644511149
transform 1 0 6440 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_66
timestamp 1644511149
transform 1 0 7176 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_70
timestamp 1644511149
transform 1 0 7544 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_77
timestamp 1644511149
transform 1 0 8188 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_83
timestamp 1644511149
transform 1 0 8740 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_84_85
timestamp 1644511149
transform 1 0 8924 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_84_91
timestamp 1644511149
transform 1 0 9476 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_116
timestamp 1644511149
transform 1 0 11776 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_84_127
timestamp 1644511149
transform 1 0 12788 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_136
timestamp 1644511149
transform 1 0 13616 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_141
timestamp 1644511149
transform 1 0 14076 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_166
timestamp 1644511149
transform 1 0 16376 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_170
timestamp 1644511149
transform 1 0 16744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_192
timestamp 1644511149
transform 1 0 18768 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_197
timestamp 1644511149
transform 1 0 19228 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_84_205
timestamp 1644511149
transform 1 0 19964 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_84_229
timestamp 1644511149
transform 1 0 22172 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_235
timestamp 1644511149
transform 1 0 22724 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_84_239
timestamp 1644511149
transform 1 0 23092 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_84_248
timestamp 1644511149
transform 1 0 23920 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_84_274
timestamp 1644511149
transform 1 0 26312 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_299
timestamp 1644511149
transform 1 0 28612 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_84_307
timestamp 1644511149
transform 1 0 29348 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_312
timestamp 1644511149
transform 1 0 29808 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_323
timestamp 1644511149
transform 1 0 30820 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_327
timestamp 1644511149
transform 1 0 31188 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_349
timestamp 1644511149
transform 1 0 33212 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_84_356
timestamp 1644511149
transform 1 0 33856 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_84_368
timestamp 1644511149
transform 1 0 34960 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_84_372
timestamp 1644511149
transform 1 0 35328 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_84_394
timestamp 1644511149
transform 1 0 37352 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_84_406
timestamp 1644511149
transform 1 0 38456 0 1 47872
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_84_418
timestamp 1644511149
transform 1 0 39560 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_84_424
timestamp 1644511149
transform 1 0 40112 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_430
timestamp 1644511149
transform 1 0 40664 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_84_434
timestamp 1644511149
transform 1 0 41032 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_84_459
timestamp 1644511149
transform 1 0 43332 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_84_469
timestamp 1644511149
transform 1 0 44252 0 1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_84_475
timestamp 1644511149
transform 1 0 44804 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_84_481
timestamp 1644511149
transform 1 0 45356 0 1 47872
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_84_489
timestamp 1644511149
transform 1 0 46092 0 1 47872
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_84_512
timestamp 1644511149
transform 1 0 48208 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_85_3
timestamp 1644511149
transform 1 0 1380 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_85_27
timestamp 1644511149
transform 1 0 3588 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_52
timestamp 1644511149
transform 1 0 5888 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_78
timestamp 1644511149
transform 1 0 8280 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_86
timestamp 1644511149
transform 1 0 9016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_108
timestamp 1644511149
transform 1 0 11040 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_116
timestamp 1644511149
transform 1 0 11776 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_85_122
timestamp 1644511149
transform 1 0 12328 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_144
timestamp 1644511149
transform 1 0 14352 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_151
timestamp 1644511149
transform 1 0 14996 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_85_159
timestamp 1644511149
transform 1 0 15732 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_164
timestamp 1644511149
transform 1 0 16192 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_190
timestamp 1644511149
transform 1 0 18584 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_197
timestamp 1644511149
transform 1 0 19228 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_85_205
timestamp 1644511149
transform 1 0 19964 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_85_211
timestamp 1644511149
transform 1 0 20516 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_220
timestamp 1644511149
transform 1 0 21344 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_228
timestamp 1644511149
transform 1 0 22080 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_253
timestamp 1644511149
transform 1 0 24380 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_260
timestamp 1644511149
transform 1 0 25024 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_269
timestamp 1644511149
transform 1 0 25852 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_276
timestamp 1644511149
transform 1 0 26496 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_281
timestamp 1644511149
transform 1 0 26956 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_303
timestamp 1644511149
transform 1 0 28980 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_85_328
timestamp 1644511149
transform 1 0 31280 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_85_358
timestamp 1644511149
transform 1 0 34040 0 -1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_85_366
timestamp 1644511149
transform 1 0 34776 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_388
timestamp 1644511149
transform 1 0 36800 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_85_393
timestamp 1644511149
transform 1 0 37260 0 -1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_85_405
timestamp 1644511149
transform 1 0 38364 0 -1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_85_410
timestamp 1644511149
transform 1 0 38824 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_85_435
timestamp 1644511149
transform 1 0 41124 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_85_444
timestamp 1644511149
transform 1 0 41952 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_449
timestamp 1644511149
transform 1 0 42412 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_453
timestamp 1644511149
transform 1 0 42780 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_475
timestamp 1644511149
transform 1 0 44804 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_85_500
timestamp 1644511149
transform 1 0 47104 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_85_505
timestamp 1644511149
transform 1 0 47564 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_85_512
timestamp 1644511149
transform 1 0 48208 0 -1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_3
timestamp 1644511149
transform 1 0 1380 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_13
timestamp 1644511149
transform 1 0 2300 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_21
timestamp 1644511149
transform 1 0 3036 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_27
timestamp 1644511149
transform 1 0 3588 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_29
timestamp 1644511149
transform 1 0 3772 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_39
timestamp 1644511149
transform 1 0 4692 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_47
timestamp 1644511149
transform 1 0 5428 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_55
timestamp 1644511149
transform 1 0 6164 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_86_57
timestamp 1644511149
transform 1 0 6348 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_80
timestamp 1644511149
transform 1 0 8464 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_106
timestamp 1644511149
transform 1 0 10856 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_86_113
timestamp 1644511149
transform 1 0 11500 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_121
timestamp 1644511149
transform 1 0 12236 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_125
timestamp 1644511149
transform 1 0 12604 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_136
timestamp 1644511149
transform 1 0 13616 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_141
timestamp 1644511149
transform 1 0 14076 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_149
timestamp 1644511149
transform 1 0 14812 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_86_156
timestamp 1644511149
transform 1 0 15456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_86_179
timestamp 1644511149
transform 1 0 17572 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_186
timestamp 1644511149
transform 1 0 18216 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_194
timestamp 1644511149
transform 1 0 18952 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_86_197
timestamp 1644511149
transform 1 0 19228 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_202
timestamp 1644511149
transform 1 0 19688 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_210
timestamp 1644511149
transform 1 0 20424 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_216
timestamp 1644511149
transform 1 0 20976 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_220
timestamp 1644511149
transform 1 0 21344 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_246
timestamp 1644511149
transform 1 0 23736 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_86_256
timestamp 1644511149
transform 1 0 24656 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_86_268
timestamp 1644511149
transform 1 0 25760 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_86_273
timestamp 1644511149
transform 1 0 26220 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_279
timestamp 1644511149
transform 1 0 26772 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_281
timestamp 1644511149
transform 1 0 26956 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_289
timestamp 1644511149
transform 1 0 27692 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_296
timestamp 1644511149
transform 1 0 28336 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_304
timestamp 1644511149
transform 1 0 29072 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_309
timestamp 1644511149
transform 1 0 29532 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_332
timestamp 1644511149
transform 1 0 31648 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_337
timestamp 1644511149
transform 1 0 32108 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_341
timestamp 1644511149
transform 1 0 32476 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_348
timestamp 1644511149
transform 1 0 33120 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_86_352
timestamp 1644511149
transform 1 0 33488 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_86_356
timestamp 1644511149
transform 1 0 33856 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_86_365
timestamp 1644511149
transform 1 0 34684 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_371
timestamp 1644511149
transform 1 0 35236 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_375
timestamp 1644511149
transform 1 0 35604 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_86_382
timestamp 1644511149
transform 1 0 36248 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_86_390
timestamp 1644511149
transform 1 0 36984 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_86_393
timestamp 1644511149
transform 1 0 37260 0 1 48960
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_86_401
timestamp 1644511149
transform 1 0 37996 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_86_406
timestamp 1644511149
transform 1 0 38456 0 1 48960
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_86_418
timestamp 1644511149
transform 1 0 39560 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_86_421
timestamp 1644511149
transform 1 0 39836 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_426
timestamp 1644511149
transform 1 0 40296 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_434
timestamp 1644511149
transform 1 0 41032 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_86_444
timestamp 1644511149
transform 1 0 41952 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_86_449
timestamp 1644511149
transform 1 0 42412 0 1 48960
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_86_472
timestamp 1644511149
transform 1 0 44528 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_86_498
timestamp 1644511149
transform 1 0 46920 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_86_505
timestamp 1644511149
transform 1 0 47564 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_86_512
timestamp 1644511149
transform 1 0 48208 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 48852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 48852 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 48852 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 48852 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 48852 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 48852 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 48852 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 48852 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 48852 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 48852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 48852 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 48852 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 48852 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 48852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 48852 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 48852 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 48852 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 48852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 48852 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 48852 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 48852 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 48852 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 48852 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 48852 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 48852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 48852 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 48852 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 48852 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 48852 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 48852 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 48852 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 48852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 48852 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 48852 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 48852 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 48852 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 48852 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 48852 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 48852 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 48852 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 48852 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 48852 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 48852 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 48852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 48852 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 48852 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 48852 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 48852 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 48852 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 48852 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 48852 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 48852 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 48852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 48852 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 48852 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 48852 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 48852 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 48852 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 48852 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 48852 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 48852 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 48852 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 48852 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 48852 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 48852 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1644511149
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1644511149
transform -1 0 48852 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1644511149
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1644511149
transform -1 0 48852 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1644511149
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1644511149
transform -1 0 48852 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1644511149
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1644511149
transform -1 0 48852 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1644511149
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1644511149
transform -1 0 48852 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1644511149
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1644511149
transform -1 0 48852 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1644511149
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1644511149
transform -1 0 48852 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1644511149
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1644511149
transform -1 0 48852 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1644511149
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1644511149
transform -1 0 48852 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1644511149
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1644511149
transform -1 0 48852 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1644511149
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1644511149
transform -1 0 48852 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1644511149
transform 1 0 1104 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1644511149
transform -1 0 48852 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1644511149
transform 1 0 1104 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1644511149
transform -1 0 48852 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_156
timestamp 1644511149
transform 1 0 1104 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_157
timestamp 1644511149
transform -1 0 48852 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_158
timestamp 1644511149
transform 1 0 1104 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_159
timestamp 1644511149
transform -1 0 48852 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_160
timestamp 1644511149
transform 1 0 1104 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_161
timestamp 1644511149
transform -1 0 48852 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_162
timestamp 1644511149
transform 1 0 1104 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_163
timestamp 1644511149
transform -1 0 48852 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_164
timestamp 1644511149
transform 1 0 1104 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_165
timestamp 1644511149
transform -1 0 48852 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_166
timestamp 1644511149
transform 1 0 1104 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_167
timestamp 1644511149
transform -1 0 48852 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_168
timestamp 1644511149
transform 1 0 1104 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_169
timestamp 1644511149
transform -1 0 48852 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_170
timestamp 1644511149
transform 1 0 1104 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_171
timestamp 1644511149
transform -1 0 48852 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_172
timestamp 1644511149
transform 1 0 1104 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_173
timestamp 1644511149
transform -1 0 48852 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 39744 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 44896 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 42320 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 47472 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 24288 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 29440 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 34592 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 39744 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 44896 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 26864 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 32016 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 37168 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 42320 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 47472 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 24288 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 29440 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 34592 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 39744 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 44896 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 26864 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 32016 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 37168 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 42320 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 47472 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 24288 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 29440 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 34592 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 39744 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 44896 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 26864 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 32016 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 37168 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 42320 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 47472 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 24288 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 29440 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 34592 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 39744 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 44896 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 26864 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 32016 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 37168 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 42320 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 47472 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_867
timestamp 1644511149
transform 1 0 3680 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_868
timestamp 1644511149
transform 1 0 8832 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_869
timestamp 1644511149
transform 1 0 13984 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_870
timestamp 1644511149
transform 1 0 19136 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_871
timestamp 1644511149
transform 1 0 24288 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_872
timestamp 1644511149
transform 1 0 29440 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_873
timestamp 1644511149
transform 1 0 34592 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_874
timestamp 1644511149
transform 1 0 39744 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_875
timestamp 1644511149
transform 1 0 44896 0 1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_876
timestamp 1644511149
transform 1 0 6256 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_877
timestamp 1644511149
transform 1 0 11408 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_878
timestamp 1644511149
transform 1 0 16560 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_879
timestamp 1644511149
transform 1 0 21712 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_880
timestamp 1644511149
transform 1 0 26864 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_881
timestamp 1644511149
transform 1 0 32016 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_882
timestamp 1644511149
transform 1 0 37168 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_883
timestamp 1644511149
transform 1 0 42320 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_884
timestamp 1644511149
transform 1 0 47472 0 -1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_885
timestamp 1644511149
transform 1 0 3680 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_886
timestamp 1644511149
transform 1 0 8832 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_887
timestamp 1644511149
transform 1 0 13984 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_888
timestamp 1644511149
transform 1 0 19136 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_889
timestamp 1644511149
transform 1 0 24288 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_890
timestamp 1644511149
transform 1 0 29440 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_891
timestamp 1644511149
transform 1 0 34592 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_892
timestamp 1644511149
transform 1 0 39744 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_893
timestamp 1644511149
transform 1 0 44896 0 1 44608
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_894
timestamp 1644511149
transform 1 0 6256 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_895
timestamp 1644511149
transform 1 0 11408 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_896
timestamp 1644511149
transform 1 0 16560 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_897
timestamp 1644511149
transform 1 0 21712 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_898
timestamp 1644511149
transform 1 0 26864 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_899
timestamp 1644511149
transform 1 0 32016 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_900
timestamp 1644511149
transform 1 0 37168 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_901
timestamp 1644511149
transform 1 0 42320 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_902
timestamp 1644511149
transform 1 0 47472 0 -1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_903
timestamp 1644511149
transform 1 0 3680 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_904
timestamp 1644511149
transform 1 0 8832 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_905
timestamp 1644511149
transform 1 0 13984 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_906
timestamp 1644511149
transform 1 0 19136 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_907
timestamp 1644511149
transform 1 0 24288 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_908
timestamp 1644511149
transform 1 0 29440 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_909
timestamp 1644511149
transform 1 0 34592 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_910
timestamp 1644511149
transform 1 0 39744 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_911
timestamp 1644511149
transform 1 0 44896 0 1 45696
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_912
timestamp 1644511149
transform 1 0 6256 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_913
timestamp 1644511149
transform 1 0 11408 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_914
timestamp 1644511149
transform 1 0 16560 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_915
timestamp 1644511149
transform 1 0 21712 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_916
timestamp 1644511149
transform 1 0 26864 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_917
timestamp 1644511149
transform 1 0 32016 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_918
timestamp 1644511149
transform 1 0 37168 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_919
timestamp 1644511149
transform 1 0 42320 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_920
timestamp 1644511149
transform 1 0 47472 0 -1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_921
timestamp 1644511149
transform 1 0 3680 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_922
timestamp 1644511149
transform 1 0 8832 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_923
timestamp 1644511149
transform 1 0 13984 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_924
timestamp 1644511149
transform 1 0 19136 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_925
timestamp 1644511149
transform 1 0 24288 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_926
timestamp 1644511149
transform 1 0 29440 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_927
timestamp 1644511149
transform 1 0 34592 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_928
timestamp 1644511149
transform 1 0 39744 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_929
timestamp 1644511149
transform 1 0 44896 0 1 46784
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_930
timestamp 1644511149
transform 1 0 6256 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_931
timestamp 1644511149
transform 1 0 11408 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_932
timestamp 1644511149
transform 1 0 16560 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_933
timestamp 1644511149
transform 1 0 21712 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_934
timestamp 1644511149
transform 1 0 26864 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_935
timestamp 1644511149
transform 1 0 32016 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_936
timestamp 1644511149
transform 1 0 37168 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_937
timestamp 1644511149
transform 1 0 42320 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_938
timestamp 1644511149
transform 1 0 47472 0 -1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_939
timestamp 1644511149
transform 1 0 3680 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_940
timestamp 1644511149
transform 1 0 8832 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_941
timestamp 1644511149
transform 1 0 13984 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_942
timestamp 1644511149
transform 1 0 19136 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_943
timestamp 1644511149
transform 1 0 24288 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_944
timestamp 1644511149
transform 1 0 29440 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_945
timestamp 1644511149
transform 1 0 34592 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_946
timestamp 1644511149
transform 1 0 39744 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_947
timestamp 1644511149
transform 1 0 44896 0 1 47872
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_948
timestamp 1644511149
transform 1 0 6256 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_949
timestamp 1644511149
transform 1 0 11408 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_950
timestamp 1644511149
transform 1 0 16560 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_951
timestamp 1644511149
transform 1 0 21712 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_952
timestamp 1644511149
transform 1 0 26864 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_953
timestamp 1644511149
transform 1 0 32016 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_954
timestamp 1644511149
transform 1 0 37168 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_955
timestamp 1644511149
transform 1 0 42320 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_956
timestamp 1644511149
transform 1 0 47472 0 -1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_957
timestamp 1644511149
transform 1 0 3680 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_958
timestamp 1644511149
transform 1 0 6256 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_959
timestamp 1644511149
transform 1 0 8832 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_960
timestamp 1644511149
transform 1 0 11408 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_961
timestamp 1644511149
transform 1 0 13984 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_962
timestamp 1644511149
transform 1 0 16560 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_963
timestamp 1644511149
transform 1 0 19136 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_964
timestamp 1644511149
transform 1 0 21712 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_965
timestamp 1644511149
transform 1 0 24288 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_966
timestamp 1644511149
transform 1 0 26864 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_967
timestamp 1644511149
transform 1 0 29440 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_968
timestamp 1644511149
transform 1 0 32016 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_969
timestamp 1644511149
transform 1 0 34592 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_970
timestamp 1644511149
transform 1 0 37168 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_971
timestamp 1644511149
transform 1 0 39744 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_972
timestamp 1644511149
transform 1 0 42320 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_973
timestamp 1644511149
transform 1 0 44896 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_974
timestamp 1644511149
transform 1 0 47472 0 1 48960
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_4  _0847_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 42432
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _0848_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_6  _0849_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27784 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__buf_12  _0850_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 1 43520
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0851_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0852_
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0853_
timestamp 1644511149
transform 1 0 2484 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0854_
timestamp 1644511149
transform 1 0 36340 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0855_
timestamp 1644511149
transform 1 0 47564 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0856_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27048 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0857_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28888 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0858_
timestamp 1644511149
transform 1 0 2208 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0859_
timestamp 1644511149
transform 1 0 43976 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0860_
timestamp 1644511149
transform 1 0 2208 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0861_
timestamp 1644511149
transform 1 0 44988 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0862_
timestamp 1644511149
transform 1 0 23644 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0863_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29900 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0864_
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0865_
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0866_
timestamp 1644511149
transform 1 0 4232 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0867_
timestamp 1644511149
transform 1 0 11592 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0868_
timestamp 1644511149
transform 1 0 45632 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0869_
timestamp 1644511149
transform 1 0 27968 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0870_
timestamp 1644511149
transform 1 0 2024 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0871_
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0872_
timestamp 1644511149
transform 1 0 22172 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0873_
timestamp 1644511149
transform 1 0 2024 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0874_
timestamp 1644511149
transform 1 0 2024 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0875_
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0876_
timestamp 1644511149
transform 1 0 37812 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0877_
timestamp 1644511149
transform 1 0 2944 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0878_
timestamp 1644511149
transform 1 0 7268 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0879_
timestamp 1644511149
transform 1 0 22540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0880_
timestamp 1644511149
transform 1 0 36524 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _0881_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27968 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0882_
timestamp 1644511149
transform 1 0 18492 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0883_
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0884_
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0885_
timestamp 1644511149
transform 1 0 30728 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0886_
timestamp 1644511149
transform 1 0 29716 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0887_
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0888_
timestamp 1644511149
transform 1 0 33580 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0889_
timestamp 1644511149
transform 1 0 33672 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0890_
timestamp 1644511149
transform 1 0 32568 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0891_
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0892_
timestamp 1644511149
transform 1 0 31004 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0893_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0894_
timestamp 1644511149
transform 1 0 32108 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0895_
timestamp 1644511149
transform 1 0 40112 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0896_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 40756 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0897_
timestamp 1644511149
transform 1 0 2668 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0898_
timestamp 1644511149
transform 1 0 2208 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0899_
timestamp 1644511149
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0900_
timestamp 1644511149
transform 1 0 31464 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0901_
timestamp 1644511149
transform 1 0 20148 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0902_
timestamp 1644511149
transform 1 0 14444 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0903_
timestamp 1644511149
transform 1 0 30176 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0904_
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0905_
timestamp 1644511149
transform 1 0 46644 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0906_
timestamp 1644511149
transform 1 0 30544 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0907_
timestamp 1644511149
transform 1 0 30544 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0908_
timestamp 1644511149
transform 1 0 2668 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0909_
timestamp 1644511149
transform 1 0 22816 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0910_
timestamp 1644511149
transform 1 0 2300 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0911_
timestamp 1644511149
transform 1 0 45632 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0912_
timestamp 1644511149
transform 1 0 29992 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0913_
timestamp 1644511149
transform 1 0 44988 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0914_
timestamp 1644511149
transform 1 0 39836 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0915_
timestamp 1644511149
transform 1 0 7268 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0916_
timestamp 1644511149
transform 1 0 46552 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0917_
timestamp 1644511149
transform 1 0 7084 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0918_
timestamp 1644511149
transform 1 0 35236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _0919_
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0920_
timestamp 1644511149
transform 1 0 33304 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0921_
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0922_
timestamp 1644511149
transform 1 0 33948 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0923_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0924_
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _0925_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 31464 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _0926_
timestamp 1644511149
transform 1 0 33580 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0927_
timestamp 1644511149
transform 1 0 33212 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0928_
timestamp 1644511149
transform 1 0 6164 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0929_
timestamp 1644511149
transform 1 0 4876 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0930_
timestamp 1644511149
transform 1 0 32384 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  _0931_
timestamp 1644511149
transform 1 0 32384 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__inv_2  _0932_
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0933_
timestamp 1644511149
transform 1 0 46828 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0934_
timestamp 1644511149
transform 1 0 2944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0935_
timestamp 1644511149
transform 1 0 41492 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0936_
timestamp 1644511149
transform 1 0 19596 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0937_
timestamp 1644511149
transform 1 0 33212 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0938_
timestamp 1644511149
transform 1 0 34684 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0939_
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0940_
timestamp 1644511149
transform 1 0 26036 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0941_
timestamp 1644511149
transform 1 0 16652 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0942_
timestamp 1644511149
transform 1 0 13340 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0943_
timestamp 1644511149
transform 1 0 32660 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0944_
timestamp 1644511149
transform 1 0 27324 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0945_
timestamp 1644511149
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0946_
timestamp 1644511149
transform 1 0 4324 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0947_
timestamp 1644511149
transform 1 0 46736 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0948_
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0949_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _0950_
timestamp 1644511149
transform 1 0 35144 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0951_
timestamp 1644511149
transform 1 0 2760 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0952_
timestamp 1644511149
transform 1 0 46644 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0953_
timestamp 1644511149
transform 1 0 46368 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0954_
timestamp 1644511149
transform 1 0 2300 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0955_
timestamp 1644511149
transform 1 0 11500 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0956_
timestamp 1644511149
transform 1 0 35972 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0957_
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0958_
timestamp 1644511149
transform 1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0959_
timestamp 1644511149
transform 1 0 37904 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0960_
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0961_
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0962_
timestamp 1644511149
transform 1 0 33396 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0963_
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0964_
timestamp 1644511149
transform 1 0 7728 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _0965_
timestamp 1644511149
transform 1 0 12880 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0966_
timestamp 1644511149
transform 1 0 45908 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0967_
timestamp 1644511149
transform 1 0 8004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _0968_
timestamp 1644511149
transform 1 0 30544 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _0969_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0970_
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0971_
timestamp 1644511149
transform 1 0 9752 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0972_
timestamp 1644511149
transform 1 0 20792 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0973_
timestamp 1644511149
transform 1 0 31004 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _0974_
timestamp 1644511149
transform 1 0 30176 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _0975_
timestamp 1644511149
transform 1 0 2944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0976_
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0977_
timestamp 1644511149
transform 1 0 8004 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0978_
timestamp 1644511149
transform 1 0 17296 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0979_
timestamp 1644511149
transform 1 0 30728 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0980_
timestamp 1644511149
transform 1 0 25300 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  _0981_
timestamp 1644511149
transform 1 0 25668 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0982_
timestamp 1644511149
transform 1 0 2944 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0983_
timestamp 1644511149
transform 1 0 28520 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0984_
timestamp 1644511149
transform 1 0 2852 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0985_
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0986_
timestamp 1644511149
transform 1 0 2208 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _0987_
timestamp 1644511149
transform 1 0 24564 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _0988_
timestamp 1644511149
transform 1 0 23276 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0989_
timestamp 1644511149
transform 1 0 23092 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0990_
timestamp 1644511149
transform 1 0 25668 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0991_
timestamp 1644511149
transform 1 0 22448 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0992_
timestamp 1644511149
transform 1 0 26220 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0993_
timestamp 1644511149
transform 1 0 26036 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _0994_
timestamp 1644511149
transform 1 0 10396 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0995_
timestamp 1644511149
transform 1 0 10212 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0996_
timestamp 1644511149
transform 1 0 11500 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0997_
timestamp 1644511149
transform 1 0 33580 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _0998_
timestamp 1644511149
transform 1 0 14260 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _0999_
timestamp 1644511149
transform 1 0 24472 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1000_
timestamp 1644511149
transform 1 0 2668 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1001_
timestamp 1644511149
transform 1 0 2024 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1002_
timestamp 1644511149
transform 1 0 2024 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1003_
timestamp 1644511149
transform 1 0 46644 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1004_
timestamp 1644511149
transform 1 0 43424 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1005_
timestamp 1644511149
transform 1 0 26036 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1006_
timestamp 1644511149
transform 1 0 2944 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1007_
timestamp 1644511149
transform 1 0 27784 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1008_
timestamp 1644511149
transform 1 0 47564 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1009_
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1010_
timestamp 1644511149
transform 1 0 46828 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1011_
timestamp 1644511149
transform 1 0 42228 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__buf_8  _1012_
timestamp 1644511149
transform 1 0 42412 0 -1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1013_
timestamp 1644511149
transform 1 0 4692 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1014_
timestamp 1644511149
transform 1 0 12512 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1015_
timestamp 1644511149
transform 1 0 26220 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1016_
timestamp 1644511149
transform 1 0 41676 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1017_
timestamp 1644511149
transform 1 0 41676 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_6  _1018_
timestamp 1644511149
transform 1 0 42412 0 -1 47872
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1019_
timestamp 1644511149
transform 1 0 3772 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1020_
timestamp 1644511149
transform 1 0 46828 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1021_
timestamp 1644511149
transform 1 0 3312 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1022_
timestamp 1644511149
transform 1 0 47564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1023_
timestamp 1644511149
transform 1 0 20148 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  _1024_
timestamp 1644511149
transform 1 0 43608 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1025_
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1026_
timestamp 1644511149
transform 1 0 45632 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1027_
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1028_
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1029_
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  _1030_
timestamp 1644511149
transform 1 0 43240 0 1 46784
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1031_
timestamp 1644511149
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1032_
timestamp 1644511149
transform 1 0 46828 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1033_
timestamp 1644511149
transform 1 0 6992 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1034_
timestamp 1644511149
transform 1 0 35788 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1035_
timestamp 1644511149
transform 1 0 47564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_12  _1036_
timestamp 1644511149
transform 1 0 41400 0 1 46784
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _1037_
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1038_
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1039_
timestamp 1644511149
transform 1 0 3772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1040_
timestamp 1644511149
transform 1 0 7912 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1041_
timestamp 1644511149
transform 1 0 29532 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1042_
timestamp 1644511149
transform 1 0 17204 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1043_
timestamp 1644511149
transform 1 0 7084 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1044_
timestamp 1644511149
transform 1 0 16836 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1045_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27232 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1046_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24840 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1047_
timestamp 1644511149
transform 1 0 23552 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1048_
timestamp 1644511149
transform 1 0 27784 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1049_
timestamp 1644511149
transform 1 0 26128 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1050_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23644 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1051_
timestamp 1644511149
transform 1 0 24748 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1052_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28796 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or4b_1  _1053_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1054_
timestamp 1644511149
transform 1 0 25484 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1055_
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1056_
timestamp 1644511149
transform 1 0 24472 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1057_
timestamp 1644511149
transform 1 0 25392 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1058_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26128 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _1059_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26220 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1060_
timestamp 1644511149
transform 1 0 14168 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1061_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1062_
timestamp 1644511149
transform 1 0 14444 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _1063_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17664 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1064_
timestamp 1644511149
transform 1 0 23828 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1065_
timestamp 1644511149
transform 1 0 29532 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1066_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18400 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _1067_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25668 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1068_
timestamp 1644511149
transform 1 0 19412 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1069_
timestamp 1644511149
transform 1 0 19412 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1070_
timestamp 1644511149
transform 1 0 17112 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1071_
timestamp 1644511149
transform 1 0 23368 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1072_
timestamp 1644511149
transform 1 0 19504 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1073_
timestamp 1644511149
transform 1 0 18952 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1074_
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a21boi_1  _1075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20056 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1076_
timestamp 1644511149
transform 1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17112 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1078_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16284 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1079_
timestamp 1644511149
transform 1 0 17020 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _1080_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1081_
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1082_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17388 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  _1083_
timestamp 1644511149
transform 1 0 25484 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1084_
timestamp 1644511149
transform 1 0 25208 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1085_
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1086_
timestamp 1644511149
transform 1 0 9292 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1087_
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1088_
timestamp 1644511149
transform 1 0 14536 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1089_
timestamp 1644511149
transform 1 0 17020 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1090_
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1091_
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1092_
timestamp 1644511149
transform 1 0 15180 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1093_
timestamp 1644511149
transform 1 0 7728 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1094_
timestamp 1644511149
transform 1 0 24380 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or4bb_2  _1095_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 47288 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or4_2  _1096_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25024 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1097_
timestamp 1644511149
transform 1 0 24656 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1098_
timestamp 1644511149
transform 1 0 24840 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _1099_
timestamp 1644511149
transform 1 0 37996 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _1100_
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1101_
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1102_
timestamp 1644511149
transform 1 0 23000 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1103_
timestamp 1644511149
transform 1 0 23460 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1104_
timestamp 1644511149
transform 1 0 23644 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1105_
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _1106_
timestamp 1644511149
transform 1 0 25300 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1107_
timestamp 1644511149
transform 1 0 19504 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1108_
timestamp 1644511149
transform 1 0 23736 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1109_
timestamp 1644511149
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and3b_4  _1110_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1111_
timestamp 1644511149
transform 1 0 18216 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1112_
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1113_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19044 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1114_
timestamp 1644511149
transform 1 0 20424 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1115_
timestamp 1644511149
transform 1 0 20240 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1116_
timestamp 1644511149
transform 1 0 20792 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1117_
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1118_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1119_
timestamp 1644511149
transform 1 0 19044 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1120_
timestamp 1644511149
transform 1 0 19412 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1121_
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1122_
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1123_
timestamp 1644511149
transform 1 0 24472 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _1124_
timestamp 1644511149
transform 1 0 20148 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1125_
timestamp 1644511149
transform 1 0 19504 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1126_
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1127_
timestamp 1644511149
transform 1 0 26128 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1128_
timestamp 1644511149
transform 1 0 27692 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1129_
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1130_
timestamp 1644511149
transform 1 0 31372 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1131_
timestamp 1644511149
transform 1 0 30268 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1132_
timestamp 1644511149
transform 1 0 31464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1133_
timestamp 1644511149
transform 1 0 30176 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1134_
timestamp 1644511149
transform 1 0 32200 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1135_
timestamp 1644511149
transform 1 0 31556 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1136_
timestamp 1644511149
transform 1 0 32384 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1137_
timestamp 1644511149
transform 1 0 26220 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1138_
timestamp 1644511149
transform 1 0 31280 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1139_
timestamp 1644511149
transform 1 0 26036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1140_
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1141_
timestamp 1644511149
transform 1 0 29348 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1142_
timestamp 1644511149
transform 1 0 29900 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1143_
timestamp 1644511149
transform 1 0 29348 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1144_
timestamp 1644511149
transform 1 0 28244 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1145_
timestamp 1644511149
transform 1 0 28428 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1146_
timestamp 1644511149
transform 1 0 27876 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1147_
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1148_
timestamp 1644511149
transform 1 0 25760 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1149_
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1150_
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1151_
timestamp 1644511149
transform 1 0 25392 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1152_
timestamp 1644511149
transform 1 0 15824 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1153_
timestamp 1644511149
transform 1 0 15732 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1154_
timestamp 1644511149
transform 1 0 18032 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1155_
timestamp 1644511149
transform 1 0 18032 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1156_
timestamp 1644511149
transform 1 0 14536 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1157_
timestamp 1644511149
transform 1 0 11960 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1158_
timestamp 1644511149
transform 1 0 12052 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1159_
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1160_
timestamp 1644511149
transform 1 0 10580 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1161_
timestamp 1644511149
transform 1 0 11960 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1162_
timestamp 1644511149
transform 1 0 17204 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1163_
timestamp 1644511149
transform 1 0 16652 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1164_
timestamp 1644511149
transform 1 0 10580 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1165_
timestamp 1644511149
transform 1 0 12236 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1166_
timestamp 1644511149
transform 1 0 11776 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1167_
timestamp 1644511149
transform 1 0 15364 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1168_
timestamp 1644511149
transform 1 0 14996 0 1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1169_
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1170_
timestamp 1644511149
transform 1 0 9292 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1171_
timestamp 1644511149
transform 1 0 8004 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1172_
timestamp 1644511149
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1173_
timestamp 1644511149
transform 1 0 7176 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1174_
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1175_
timestamp 1644511149
transform 1 0 9200 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1176_
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1177_
timestamp 1644511149
transform 1 0 14168 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1178_
timestamp 1644511149
transform 1 0 23552 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1179_
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1180_
timestamp 1644511149
transform 1 0 14996 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or4_1  _1181_
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1182_
timestamp 1644511149
transform 1 0 20976 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1183_
timestamp 1644511149
transform 1 0 16284 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1184_
timestamp 1644511149
transform 1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1185_
timestamp 1644511149
transform 1 0 16744 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1186_
timestamp 1644511149
transform 1 0 14260 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1187_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1188_
timestamp 1644511149
transform 1 0 19504 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1189_
timestamp 1644511149
transform 1 0 13156 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1190_
timestamp 1644511149
transform 1 0 13432 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1191_
timestamp 1644511149
transform 1 0 14076 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1192_
timestamp 1644511149
transform 1 0 14444 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1193_
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1194_
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1195_
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1196_
timestamp 1644511149
transform 1 0 17756 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1197_
timestamp 1644511149
transform 1 0 13340 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1198_
timestamp 1644511149
transform 1 0 16652 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1199_
timestamp 1644511149
transform 1 0 19780 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1200_
timestamp 1644511149
transform 1 0 19228 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1201_
timestamp 1644511149
transform 1 0 20148 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1202_
timestamp 1644511149
transform 1 0 20332 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1203_
timestamp 1644511149
transform 1 0 17664 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1204_
timestamp 1644511149
transform 1 0 17848 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1205_
timestamp 1644511149
transform 1 0 16376 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1206_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1207_
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1208_
timestamp 1644511149
transform 1 0 20424 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1209_
timestamp 1644511149
transform 1 0 20516 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1210_
timestamp 1644511149
transform 1 0 22448 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1211_
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _1212_
timestamp 1644511149
transform 1 0 21068 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1213_
timestamp 1644511149
transform 1 0 22172 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1214_
timestamp 1644511149
transform 1 0 21988 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1215_
timestamp 1644511149
transform 1 0 19964 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1216_
timestamp 1644511149
transform 1 0 23092 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1217_
timestamp 1644511149
transform 1 0 23184 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1218_
timestamp 1644511149
transform 1 0 20424 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _1219_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19412 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1220_
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1221_
timestamp 1644511149
transform 1 0 20884 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1222_
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1223_
timestamp 1644511149
transform 1 0 23184 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1224_
timestamp 1644511149
transform 1 0 28612 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1225_
timestamp 1644511149
transform 1 0 27876 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1226_
timestamp 1644511149
transform 1 0 28612 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1227_
timestamp 1644511149
transform 1 0 20608 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1228_
timestamp 1644511149
transform 1 0 23920 0 -1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1229_
timestamp 1644511149
transform 1 0 33580 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1230_
timestamp 1644511149
transform 1 0 33488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1231_
timestamp 1644511149
transform 1 0 32660 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1232_
timestamp 1644511149
transform 1 0 33764 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1233_
timestamp 1644511149
transform 1 0 33672 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1234_
timestamp 1644511149
transform 1 0 33948 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1235_
timestamp 1644511149
transform 1 0 30176 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1236_
timestamp 1644511149
transform 1 0 29072 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1237_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1238_
timestamp 1644511149
transform 1 0 19596 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1239_
timestamp 1644511149
transform 1 0 21344 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1240_
timestamp 1644511149
transform 1 0 18952 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1241_
timestamp 1644511149
transform 1 0 18032 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1242_
timestamp 1644511149
transform 1 0 19136 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1243_
timestamp 1644511149
transform 1 0 18032 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1244_
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1245_
timestamp 1644511149
transform 1 0 17940 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1246_
timestamp 1644511149
transform 1 0 19780 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1247_
timestamp 1644511149
transform 1 0 20240 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1248_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23920 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _1249_
timestamp 1644511149
transform 1 0 7636 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1250_
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1251_
timestamp 1644511149
transform 1 0 24564 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1252_
timestamp 1644511149
transform 1 0 24748 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1253_
timestamp 1644511149
transform 1 0 28704 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_2  _1254_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1255_
timestamp 1644511149
transform 1 0 27784 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1256_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2b_1  _1257_
timestamp 1644511149
transform 1 0 24012 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o221a_1  _1258_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23092 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1259_
timestamp 1644511149
transform 1 0 26956 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1260_
timestamp 1644511149
transform 1 0 23644 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1261_
timestamp 1644511149
transform 1 0 23644 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1262_
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1263_
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1264_
timestamp 1644511149
transform 1 0 25024 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1265_
timestamp 1644511149
transform 1 0 25208 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1266_
timestamp 1644511149
transform 1 0 24012 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1267_
timestamp 1644511149
transform 1 0 23276 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1268_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23276 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1269_
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1270_
timestamp 1644511149
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1271_
timestamp 1644511149
transform 1 0 24840 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o22a_1  _1272_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22632 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1273_
timestamp 1644511149
transform 1 0 22448 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1274_
timestamp 1644511149
transform 1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1275_
timestamp 1644511149
transform 1 0 27784 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1276_
timestamp 1644511149
transform 1 0 25668 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1277_
timestamp 1644511149
transform 1 0 24656 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1278_
timestamp 1644511149
transform 1 0 27968 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1279_
timestamp 1644511149
transform 1 0 25208 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1280_
timestamp 1644511149
transform 1 0 30912 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1281_
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1282_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25760 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1283_
timestamp 1644511149
transform 1 0 26036 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1284_
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1285_
timestamp 1644511149
transform 1 0 26128 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1286_
timestamp 1644511149
transform 1 0 25668 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _1287_
timestamp 1644511149
transform 1 0 28704 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1288_
timestamp 1644511149
transform 1 0 27968 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1289_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28428 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1290_
timestamp 1644511149
transform 1 0 27600 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1291_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28336 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1292_
timestamp 1644511149
transform 1 0 28152 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1293_
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1294_
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1295_
timestamp 1644511149
transform 1 0 28244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1296_
timestamp 1644511149
transform 1 0 29440 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1297_
timestamp 1644511149
transform 1 0 29716 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1298_
timestamp 1644511149
transform 1 0 30176 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__or4_2  _1299_
timestamp 1644511149
transform 1 0 28980 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1300_
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1301_
timestamp 1644511149
transform 1 0 29532 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1302_
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1303_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1304_
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__and2b_1  _1305_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30084 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1306_
timestamp 1644511149
transform 1 0 30452 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1307_
timestamp 1644511149
transform 1 0 31004 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1308_
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1309_
timestamp 1644511149
transform 1 0 32844 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _1310_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 30636 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1311_
timestamp 1644511149
transform 1 0 31188 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1312_
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1313_
timestamp 1644511149
transform 1 0 29808 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1314_
timestamp 1644511149
transform 1 0 30820 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1315_
timestamp 1644511149
transform 1 0 30452 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1316_
timestamp 1644511149
transform 1 0 30360 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _1317_
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1318_
timestamp 1644511149
transform 1 0 29440 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o221a_1  _1319_
timestamp 1644511149
transform 1 0 32752 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1320_
timestamp 1644511149
transform 1 0 29624 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1321_
timestamp 1644511149
transform 1 0 28612 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _1322_
timestamp 1644511149
transform 1 0 29348 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1323_
timestamp 1644511149
transform 1 0 27416 0 -1 17408
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _1324_
timestamp 1644511149
transform 1 0 28520 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1325_
timestamp 1644511149
transform 1 0 28704 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1326_
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1327_
timestamp 1644511149
transform 1 0 29808 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1328_
timestamp 1644511149
transform 1 0 27232 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1329_
timestamp 1644511149
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1330_
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _1331_
timestamp 1644511149
transform 1 0 27508 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1332_
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o21a_1  _1333_
timestamp 1644511149
transform 1 0 25668 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1334_
timestamp 1644511149
transform 1 0 24748 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1335_
timestamp 1644511149
transform 1 0 25300 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_1  _1336_
timestamp 1644511149
transform 1 0 25944 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1337_
timestamp 1644511149
transform 1 0 24748 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1338_
timestamp 1644511149
transform 1 0 26036 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1339_
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1340_
timestamp 1644511149
transform 1 0 23644 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1341_
timestamp 1644511149
transform 1 0 22448 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1342_
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1343_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1344_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22540 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1345_
timestamp 1644511149
transform 1 0 22172 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1346_
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1347_
timestamp 1644511149
transform 1 0 23368 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _1348_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21620 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1349_
timestamp 1644511149
transform 1 0 22908 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1350_
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1351_
timestamp 1644511149
transform 1 0 22080 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1352_
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1353_
timestamp 1644511149
transform 1 0 24840 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1354_
timestamp 1644511149
transform 1 0 23092 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1355_
timestamp 1644511149
transform 1 0 25484 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1356_
timestamp 1644511149
transform 1 0 24932 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1357_
timestamp 1644511149
transform 1 0 23736 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _1358_
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _1359_
timestamp 1644511149
transform 1 0 25852 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1360_
timestamp 1644511149
transform 1 0 25852 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__or4_1  _1361_
timestamp 1644511149
transform 1 0 24748 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1362_
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1363_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 25300 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1364_
timestamp 1644511149
transform 1 0 26128 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1365_
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1366_
timestamp 1644511149
transform 1 0 25392 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1367_
timestamp 1644511149
transform 1 0 24472 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1368_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1369_
timestamp 1644511149
transform 1 0 25208 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or4_2  _1370_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1371_
timestamp 1644511149
transform 1 0 9292 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1372_
timestamp 1644511149
transform 1 0 9660 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _1373_
timestamp 1644511149
transform 1 0 9660 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_1  _1374_
timestamp 1644511149
transform 1 0 9200 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3b_1  _1375_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7912 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1376_
timestamp 1644511149
transform 1 0 7544 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1377_
timestamp 1644511149
transform 1 0 9016 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211oi_1  _1378_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1379_
timestamp 1644511149
transform 1 0 9292 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1380_
timestamp 1644511149
transform 1 0 10304 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1381_
timestamp 1644511149
transform 1 0 10396 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1382_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1383_
timestamp 1644511149
transform 1 0 14076 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1384_
timestamp 1644511149
transform 1 0 12696 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _1385_
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1386_
timestamp 1644511149
transform 1 0 12512 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _1387_
timestamp 1644511149
transform 1 0 10120 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1388_
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1389_
timestamp 1644511149
transform 1 0 13340 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1390_
timestamp 1644511149
transform 1 0 14076 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1391_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1392_
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1393_
timestamp 1644511149
transform 1 0 13248 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1394_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1395_
timestamp 1644511149
transform 1 0 13432 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__or4_1  _1396_
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _1397_
timestamp 1644511149
transform 1 0 12512 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1398_
timestamp 1644511149
transform 1 0 13064 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_1  _1399_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11776 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1400_
timestamp 1644511149
transform 1 0 11592 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _1401_
timestamp 1644511149
transform 1 0 15548 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1402_
timestamp 1644511149
transform 1 0 14812 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2b_1  _1403_
timestamp 1644511149
transform 1 0 14352 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1404_
timestamp 1644511149
transform 1 0 12880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1405_
timestamp 1644511149
transform 1 0 11500 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1406_
timestamp 1644511149
transform 1 0 13984 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1407_
timestamp 1644511149
transform 1 0 14260 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1408_
timestamp 1644511149
transform 1 0 13524 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1409_
timestamp 1644511149
transform 1 0 23552 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _1410_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 13064 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1411_
timestamp 1644511149
transform 1 0 12972 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1412_
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1413_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand3_1  _1414_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15180 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1415_
timestamp 1644511149
transform 1 0 14260 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o2111a_1  _1416_
timestamp 1644511149
transform 1 0 13064 0 -1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1417_
timestamp 1644511149
transform 1 0 13156 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1418_
timestamp 1644511149
transform 1 0 12972 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1419_
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o2111a_1  _1420_
timestamp 1644511149
transform 1 0 11776 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1421_
timestamp 1644511149
transform 1 0 10120 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1422_
timestamp 1644511149
transform 1 0 10764 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1423_
timestamp 1644511149
transform 1 0 10580 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _1424_
timestamp 1644511149
transform 1 0 10488 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1425_
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1426_
timestamp 1644511149
transform 1 0 9844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1427_
timestamp 1644511149
transform 1 0 10856 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1428_
timestamp 1644511149
transform 1 0 10212 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1429_
timestamp 1644511149
transform 1 0 9476 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o2111a_1  _1430_
timestamp 1644511149
transform 1 0 10304 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _1431_
timestamp 1644511149
transform 1 0 9844 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1432_
timestamp 1644511149
transform 1 0 10856 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1433_
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1434_
timestamp 1644511149
transform 1 0 18492 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1435_
timestamp 1644511149
transform 1 0 25760 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1436_
timestamp 1644511149
transform 1 0 19596 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1437_
timestamp 1644511149
transform 1 0 26128 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__mux2_1  _1438_
timestamp 1644511149
transform 1 0 27600 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1439_
timestamp 1644511149
transform 1 0 25484 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1440_
timestamp 1644511149
transform 1 0 25576 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1441_
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1442_
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1443_
timestamp 1644511149
transform 1 0 28612 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1444_
timestamp 1644511149
transform 1 0 28612 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1445_
timestamp 1644511149
transform 1 0 25024 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1446_
timestamp 1644511149
transform 1 0 28336 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1447_
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1448_
timestamp 1644511149
transform 1 0 27784 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1449_
timestamp 1644511149
transform 1 0 29072 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1450_
timestamp 1644511149
transform 1 0 28520 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1451_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1452_
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1453_
timestamp 1644511149
transform 1 0 29164 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1454_
timestamp 1644511149
transform 1 0 28336 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1455_
timestamp 1644511149
transform 1 0 29716 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1456_
timestamp 1644511149
transform 1 0 19596 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1457_
timestamp 1644511149
transform 1 0 28060 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1458_
timestamp 1644511149
transform 1 0 27232 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1459_
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1460_
timestamp 1644511149
transform 1 0 20608 0 1 31552
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1461_
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1462_
timestamp 1644511149
transform 1 0 24380 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1463_
timestamp 1644511149
transform 1 0 23000 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1464_
timestamp 1644511149
transform 1 0 24748 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1465_
timestamp 1644511149
transform 1 0 22816 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1466_
timestamp 1644511149
transform 1 0 21620 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1467_
timestamp 1644511149
transform 1 0 20884 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1468_
timestamp 1644511149
transform 1 0 20332 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1469_
timestamp 1644511149
transform 1 0 20700 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1470_
timestamp 1644511149
transform 1 0 20332 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1471_
timestamp 1644511149
transform 1 0 19596 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1472_
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1473_
timestamp 1644511149
transform 1 0 23460 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1474_
timestamp 1644511149
transform 1 0 25116 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1475_
timestamp 1644511149
transform 1 0 18400 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1476_
timestamp 1644511149
transform 1 0 22264 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1644511149
transform 1 0 21896 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1478_
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1479_
timestamp 1644511149
transform 1 0 23644 0 -1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1480_
timestamp 1644511149
transform 1 0 27876 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1481_
timestamp 1644511149
transform 1 0 24932 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1482_
timestamp 1644511149
transform 1 0 23460 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1483_
timestamp 1644511149
transform 1 0 22172 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1484_
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1485_
timestamp 1644511149
transform 1 0 25300 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1486_
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1487_
timestamp 1644511149
transform 1 0 26864 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1488_
timestamp 1644511149
transform 1 0 25576 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1489_
timestamp 1644511149
transform 1 0 24748 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1490_
timestamp 1644511149
transform 1 0 26772 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1491_
timestamp 1644511149
transform 1 0 24288 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 1644511149
transform 1 0 23460 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1493_
timestamp 1644511149
transform 1 0 21988 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1494_
timestamp 1644511149
transform 1 0 16928 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1495_
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1496_
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1497_
timestamp 1644511149
transform 1 0 20608 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1498_
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1499_
timestamp 1644511149
transform 1 0 23460 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1500_
timestamp 1644511149
transform 1 0 19228 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1501_
timestamp 1644511149
transform 1 0 19228 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1502_
timestamp 1644511149
transform 1 0 21344 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _1503_
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1504_
timestamp 1644511149
transform 1 0 22540 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1505_
timestamp 1644511149
transform 1 0 20424 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1506_
timestamp 1644511149
transform 1 0 21252 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1507_
timestamp 1644511149
transform 1 0 21620 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1508_
timestamp 1644511149
transform 1 0 20792 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1509_
timestamp 1644511149
transform 1 0 20608 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1510_
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1511_
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1512_
timestamp 1644511149
transform 1 0 17664 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1513_
timestamp 1644511149
transform 1 0 18216 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1514_
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1515_
timestamp 1644511149
transform 1 0 18216 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1516_
timestamp 1644511149
transform 1 0 17664 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1517_
timestamp 1644511149
transform 1 0 24380 0 1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1518_
timestamp 1644511149
transform 1 0 24012 0 -1 39168
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1519_
timestamp 1644511149
transform 1 0 22724 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1520_
timestamp 1644511149
transform 1 0 24564 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1521_
timestamp 1644511149
transform 1 0 27324 0 -1 39168
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1522_
timestamp 1644511149
transform 1 0 27508 0 1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1523_
timestamp 1644511149
transform 1 0 28336 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _1524_
timestamp 1644511149
transform 1 0 26956 0 -1 40256
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 1644511149
transform 1 0 28152 0 -1 40256
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1526_
timestamp 1644511149
transform 1 0 28336 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1644511149
transform 1 0 29624 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1528_
timestamp 1644511149
transform 1 0 28888 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1529_
timestamp 1644511149
transform 1 0 18308 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1530_
timestamp 1644511149
transform 1 0 20516 0 1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__a21o_1  _1531_
timestamp 1644511149
transform 1 0 22540 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1532_
timestamp 1644511149
transform 1 0 22632 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1533_
timestamp 1644511149
transform 1 0 21620 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1534_
timestamp 1644511149
transform 1 0 19596 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1535_
timestamp 1644511149
transform 1 0 21804 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1536_
timestamp 1644511149
transform 1 0 19412 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1537_
timestamp 1644511149
transform 1 0 19228 0 1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1538_
timestamp 1644511149
transform 1 0 19964 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1539_
timestamp 1644511149
transform 1 0 18860 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1540_
timestamp 1644511149
transform 1 0 22540 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1541_
timestamp 1644511149
transform 1 0 23092 0 1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1542_
timestamp 1644511149
transform 1 0 25668 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1543_
timestamp 1644511149
transform 1 0 25668 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1544_
timestamp 1644511149
transform 1 0 19412 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1545_
timestamp 1644511149
transform 1 0 17480 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1546_
timestamp 1644511149
transform 1 0 17388 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1547_
timestamp 1644511149
transform 1 0 27692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1548_
timestamp 1644511149
transform 1 0 27324 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1549_
timestamp 1644511149
transform 1 0 29900 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1644511149
transform 1 0 27968 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1551_
timestamp 1644511149
transform 1 0 27324 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1552_
timestamp 1644511149
transform 1 0 31188 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1553_
timestamp 1644511149
transform 1 0 31372 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1644511149
transform 1 0 32200 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1555_
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1556_
timestamp 1644511149
transform 1 0 29164 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1557_
timestamp 1644511149
transform 1 0 28980 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1558_
timestamp 1644511149
transform 1 0 32200 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1559_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1560_
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1561_
timestamp 1644511149
transform 1 0 30912 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1562_
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1563_
timestamp 1644511149
transform 1 0 30636 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1564_
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1565_
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1566_
timestamp 1644511149
transform 1 0 17020 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1567_
timestamp 1644511149
transform 1 0 15732 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__or2_1  _1568_
timestamp 1644511149
transform 1 0 16652 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1569_
timestamp 1644511149
transform 1 0 15456 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1570_
timestamp 1644511149
transform 1 0 18860 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1571_
timestamp 1644511149
transform 1 0 18032 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1572_
timestamp 1644511149
transform 1 0 17480 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1573_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1644511149
transform 1 0 19044 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1575_
timestamp 1644511149
transform 1 0 17940 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1576_
timestamp 1644511149
transform 1 0 19688 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1577_
timestamp 1644511149
transform 1 0 19596 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_1  _1578_
timestamp 1644511149
transform 1 0 18032 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1579_
timestamp 1644511149
transform 1 0 15824 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1580_
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1581_
timestamp 1644511149
transform 1 0 8004 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1582_
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1644511149
transform 1 0 8096 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1584_
timestamp 1644511149
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1585_
timestamp 1644511149
transform 1 0 17480 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1586_
timestamp 1644511149
transform 1 0 17572 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1587_
timestamp 1644511149
transform 1 0 17480 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__dfxtp_1  _1588_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 21528 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1589_
timestamp 1644511149
transform 1 0 16744 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1590_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1591_
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1592_
timestamp 1644511149
transform 1 0 17296 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1593_
timestamp 1644511149
transform 1 0 20608 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1594_
timestamp 1644511149
transform 1 0 19780 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1595_
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1596_
timestamp 1644511149
transform 1 0 17296 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1597_
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1598_
timestamp 1644511149
transform 1 0 30176 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1599_
timestamp 1644511149
transform 1 0 29624 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1600_
timestamp 1644511149
transform 1 0 32200 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1601_
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1602_
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1603_
timestamp 1644511149
transform 1 0 27600 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1604_
timestamp 1644511149
transform 1 0 27600 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1605_
timestamp 1644511149
transform 1 0 25760 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1606_
timestamp 1644511149
transform 1 0 25576 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1607_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1608_
timestamp 1644511149
transform 1 0 10396 0 1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1609_
timestamp 1644511149
transform 1 0 10120 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1610_
timestamp 1644511149
transform 1 0 16744 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1611_
timestamp 1644511149
transform 1 0 10672 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1612_
timestamp 1644511149
transform 1 0 7452 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1613_
timestamp 1644511149
transform 1 0 7820 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1614_
timestamp 1644511149
transform 1 0 7820 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1615_
timestamp 1644511149
transform 1 0 7360 0 -1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1616_
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1617_
timestamp 1644511149
transform 1 0 15364 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1618_
timestamp 1644511149
transform 1 0 13156 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1619_
timestamp 1644511149
transform 1 0 14260 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1620_
timestamp 1644511149
transform 1 0 16100 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1621_
timestamp 1644511149
transform 1 0 13156 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1622_
timestamp 1644511149
transform 1 0 19688 0 1 23936
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1623_
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1624_
timestamp 1644511149
transform 1 0 15548 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1625_
timestamp 1644511149
transform 1 0 20516 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1626_
timestamp 1644511149
transform 1 0 21804 0 -1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1627_
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1628_
timestamp 1644511149
transform 1 0 23644 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1629_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1630_
timestamp 1644511149
transform 1 0 21068 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1631_
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1632_
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1633_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1634_
timestamp 1644511149
transform 1 0 33764 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1635_
timestamp 1644511149
transform 1 0 34684 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1636_
timestamp 1644511149
transform 1 0 30176 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1637_
timestamp 1644511149
transform 1 0 22080 0 -1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1638_
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1639_
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1640_
timestamp 1644511149
transform 1 0 18032 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1641_
timestamp 1644511149
transform 1 0 21160 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1642_
timestamp 1644511149
transform 1 0 6808 0 1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1643_
timestamp 1644511149
transform 1 0 23092 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1644_
timestamp 1644511149
transform 1 0 22172 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1645_
timestamp 1644511149
transform 1 0 21344 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1646_
timestamp 1644511149
transform 1 0 26128 0 1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1647_
timestamp 1644511149
transform 1 0 25944 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1648_
timestamp 1644511149
transform 1 0 28336 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1649_
timestamp 1644511149
transform 1 0 30544 0 1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1650_
timestamp 1644511149
transform 1 0 30728 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1651_
timestamp 1644511149
transform 1 0 32384 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1652_
timestamp 1644511149
transform 1 0 32568 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1653_
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1654_
timestamp 1644511149
transform 1 0 30912 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1655_
timestamp 1644511149
transform 1 0 27600 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1656_
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1657_
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1658_
timestamp 1644511149
transform 1 0 21068 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1659_
timestamp 1644511149
transform 1 0 15364 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1660_
timestamp 1644511149
transform 1 0 25024 0 -1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1661_
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1662_
timestamp 1644511149
transform 1 0 14168 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1663_
timestamp 1644511149
transform 1 0 12696 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1664_
timestamp 1644511149
transform 1 0 11592 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1665_
timestamp 1644511149
transform 1 0 9568 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1666_
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1667_
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1668_
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1669_
timestamp 1644511149
transform 1 0 25760 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1670_
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1671_
timestamp 1644511149
transform 1 0 30084 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1672_
timestamp 1644511149
transform 1 0 28612 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1673_
timestamp 1644511149
transform 1 0 30360 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1674_
timestamp 1644511149
transform 1 0 26956 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1675_
timestamp 1644511149
transform 1 0 22908 0 -1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1676_
timestamp 1644511149
transform 1 0 20700 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1677_
timestamp 1644511149
transform 1 0 19596 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1678_
timestamp 1644511149
transform 1 0 25760 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1679_
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1680_
timestamp 1644511149
transform 1 0 23920 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1681_
timestamp 1644511149
transform 1 0 27784 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1682_
timestamp 1644511149
transform 1 0 27324 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1683_
timestamp 1644511149
transform 1 0 22448 0 -1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1684_
timestamp 1644511149
transform 1 0 20976 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1685_
timestamp 1644511149
transform 1 0 17848 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1686_
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1687_
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1688_
timestamp 1644511149
transform 1 0 17756 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1689_
timestamp 1644511149
transform 1 0 17296 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1690_
timestamp 1644511149
transform 1 0 24472 0 1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1691_
timestamp 1644511149
transform 1 0 29532 0 1 38080
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1692_
timestamp 1644511149
transform 1 0 28520 0 -1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1693_
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1694_
timestamp 1644511149
transform 1 0 22724 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1695_
timestamp 1644511149
transform 1 0 21252 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1696_
timestamp 1644511149
transform 1 0 19044 0 -1 40256
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1697_
timestamp 1644511149
transform 1 0 19228 0 1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1698_
timestamp 1644511149
transform 1 0 23184 0 -1 41344
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1699_
timestamp 1644511149
transform 1 0 26220 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1700_
timestamp 1644511149
transform 1 0 17296 0 1 39168
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_2  _1701_
timestamp 1644511149
transform 1 0 27232 0 1 27200
box -38 -48 1602 592
use sky130_fd_sc_hd__dfxtp_1  _1702_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1703_
timestamp 1644511149
transform 1 0 32476 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1704_
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1705_
timestamp 1644511149
transform 1 0 32476 0 1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1706_
timestamp 1644511149
transform 1 0 31740 0 1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1707_
timestamp 1644511149
transform 1 0 32200 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1708_
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1709_
timestamp 1644511149
transform 1 0 14904 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1710_
timestamp 1644511149
transform 1 0 19044 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1711_
timestamp 1644511149
transform 1 0 16376 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1712_
timestamp 1644511149
transform 1 0 19688 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1713_
timestamp 1644511149
transform 1 0 19412 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1714_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1715_
timestamp 1644511149
transform 1 0 7084 0 -1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1716_
timestamp 1644511149
transform 1 0 6808 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_4  _1717_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18124 0 -1 30464
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxtp_1  _1718_
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1719_
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  _1720_
timestamp 1644511149
transform 1 0 16192 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__conb_1  _1721__200 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 39928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1722__201
timestamp 1644511149
transform 1 0 32200 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1723__202
timestamp 1644511149
transform 1 0 9200 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1724__203
timestamp 1644511149
transform 1 0 1840 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1725__96
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1726__97
timestamp 1644511149
transform 1 0 26220 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1727__98
timestamp 1644511149
transform 1 0 15916 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1728__99
timestamp 1644511149
transform 1 0 25760 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1729__100
timestamp 1644511149
transform 1 0 35328 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1730__101
timestamp 1644511149
transform 1 0 2116 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1731__102
timestamp 1644511149
transform 1 0 46828 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1732__103
timestamp 1644511149
transform 1 0 1472 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1733__104
timestamp 1644511149
transform 1 0 1840 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1734__105
timestamp 1644511149
transform 1 0 2668 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1735__106
timestamp 1644511149
transform 1 0 30912 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1736__107
timestamp 1644511149
transform 1 0 17940 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1737__108
timestamp 1644511149
transform 1 0 2668 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1738__109
timestamp 1644511149
transform 1 0 32844 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1739__110
timestamp 1644511149
transform 1 0 5244 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1740__111
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1741__112
timestamp 1644511149
transform 1 0 23460 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1742__113
timestamp 1644511149
transform 1 0 12512 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1743__114
timestamp 1644511149
transform 1 0 29808 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1744__115
timestamp 1644511149
transform 1 0 20240 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1745__116
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1746__117
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1747__118
timestamp 1644511149
transform 1 0 5336 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1748__119
timestamp 1644511149
transform 1 0 40756 0 1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1749__120
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1750__121
timestamp 1644511149
transform 1 0 1564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1751__122
timestamp 1644511149
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1752__123
timestamp 1644511149
transform 1 0 20240 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1753__124
timestamp 1644511149
transform 1 0 15088 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1754__125
timestamp 1644511149
transform 1 0 30268 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1755__126
timestamp 1644511149
transform 1 0 2852 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1756__127
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1757__128
timestamp 1644511149
transform 1 0 30268 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1758__129
timestamp 1644511149
transform 1 0 2484 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1759__130
timestamp 1644511149
transform 1 0 21804 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1760__131
timestamp 1644511149
transform 1 0 1656 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1761__132
timestamp 1644511149
transform 1 0 47196 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1762__133
timestamp 1644511149
transform 1 0 1380 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1763__134
timestamp 1644511149
transform 1 0 47564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1764__135
timestamp 1644511149
transform 1 0 44252 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1765__136
timestamp 1644511149
transform 1 0 46828 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1766__137
timestamp 1644511149
transform 1 0 3404 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1767__138
timestamp 1644511149
transform 1 0 35972 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1768__139
timestamp 1644511149
transform 1 0 12512 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1769__140
timestamp 1644511149
transform 1 0 46828 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1770__141
timestamp 1644511149
transform 1 0 44252 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1771__142
timestamp 1644511149
transform 1 0 38548 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1772__143
timestamp 1644511149
transform 1 0 11500 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1773__144
timestamp 1644511149
transform 1 0 6808 0 1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1774__145
timestamp 1644511149
transform 1 0 46184 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1775__146
timestamp 1644511149
transform 1 0 33580 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1776__147
timestamp 1644511149
transform 1 0 14720 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1777__148
timestamp 1644511149
transform 1 0 2944 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1778__149
timestamp 1644511149
transform 1 0 1840 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1779__150
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1780__151
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1781__152
timestamp 1644511149
transform 1 0 43608 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1782__153
timestamp 1644511149
transform 1 0 2116 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1783__154
timestamp 1644511149
transform 1 0 28060 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1784__155
timestamp 1644511149
transform 1 0 46184 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1785__156
timestamp 1644511149
transform 1 0 42872 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1786__157
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1787__158
timestamp 1644511149
transform 1 0 4048 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1788__159
timestamp 1644511149
transform 1 0 13156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1789__160
timestamp 1644511149
transform 1 0 25576 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1790__161
timestamp 1644511149
transform 1 0 41032 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1791__162
timestamp 1644511149
transform 1 0 6072 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1792__163
timestamp 1644511149
transform 1 0 40020 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1793__164
timestamp 1644511149
transform 1 0 5152 0 -1 46784
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1794__165
timestamp 1644511149
transform 1 0 46552 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1795__166
timestamp 1644511149
transform 1 0 2668 0 1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1796__167
timestamp 1644511149
transform 1 0 46828 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1797__168
timestamp 1644511149
transform 1 0 20792 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1798__169
timestamp 1644511149
transform 1 0 47472 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1799__170
timestamp 1644511149
transform 1 0 44528 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1800__171
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1801__172
timestamp 1644511149
transform 1 0 46828 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1802__173
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1803__174
timestamp 1644511149
transform 1 0 6716 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1804__175
timestamp 1644511149
transform 1 0 45632 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1805__176
timestamp 1644511149
transform 1 0 8648 0 -1 47872
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1806__177
timestamp 1644511149
transform 1 0 46828 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1807__178
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1808__179
timestamp 1644511149
transform 1 0 1840 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1809__180
timestamp 1644511149
transform 1 0 1840 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1810__181
timestamp 1644511149
transform 1 0 36064 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1811__182
timestamp 1644511149
transform 1 0 44988 0 1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1812__183
timestamp 1644511149
transform 1 0 3312 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1813__184
timestamp 1644511149
transform 1 0 43608 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1814__185
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1815__186
timestamp 1644511149
transform 1 0 45080 0 -1 44608
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1816__187
timestamp 1644511149
transform 1 0 24748 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1817__188
timestamp 1644511149
transform 1 0 1840 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1818__189
timestamp 1644511149
transform 1 0 46828 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1819__190
timestamp 1644511149
transform 1 0 3772 0 1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1820__191
timestamp 1644511149
transform 1 0 11776 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1821__192
timestamp 1644511149
transform 1 0 43884 0 -1 45696
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1822__193
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1823__194
timestamp 1644511149
transform 1 0 32200 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1824__195
timestamp 1644511149
transform 1 0 21068 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1825__196
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1826__197
timestamp 1644511149
transform 1 0 1840 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1827__198
timestamp 1644511149
transform 1 0 38548 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  _1828__199
timestamp 1644511149
transform 1 0 2116 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__ebufn_8  _1829_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1830_
timestamp 1644511149
transform 1 0 16744 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1831_
timestamp 1644511149
transform 1 0 21988 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1832_
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1833_
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1834_
timestamp 1644511149
transform 1 0 18860 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1835_
timestamp 1644511149
transform 1 0 26496 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1836_
timestamp 1644511149
transform 1 0 31372 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1837_
timestamp 1644511149
transform 1 0 29624 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1838_
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1839_
timestamp 1644511149
transform 1 0 32752 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1840_
timestamp 1644511149
transform 1 0 32844 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1841_
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1842_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1843_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1844_
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1845_
timestamp 1644511149
transform 1 0 20332 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1846_
timestamp 1644511149
transform 1 0 7728 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1847_
timestamp 1644511149
transform 1 0 10396 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1848_
timestamp 1644511149
transform 1 0 23000 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1849_
timestamp 1644511149
transform 1 0 10948 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1850_
timestamp 1644511149
transform 1 0 2668 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1851_
timestamp 1644511149
transform 1 0 7912 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1852_
timestamp 1644511149
transform 1 0 3680 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1853_
timestamp 1644511149
transform 1 0 6256 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1854_
timestamp 1644511149
transform 1 0 10580 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1855_
timestamp 1644511149
transform 1 0 3496 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1856_
timestamp 1644511149
transform 1 0 27048 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1857_
timestamp 1644511149
transform 1 0 16652 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1858_
timestamp 1644511149
transform 1 0 25668 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1859_
timestamp 1644511149
transform 1 0 34868 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1860_
timestamp 1644511149
transform 1 0 2024 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1861_
timestamp 1644511149
transform 1 0 46276 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_2  _1862_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6624 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__ebufn_8  _1863_
timestamp 1644511149
transform 1 0 17112 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1864_
timestamp 1644511149
transform 1 0 29348 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1865_
timestamp 1644511149
transform 1 0 6348 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1866_
timestamp 1644511149
transform 1 0 1380 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1867_
timestamp 1644511149
transform 1 0 40572 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1868_
timestamp 1644511149
transform 1 0 32108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1869_
timestamp 1644511149
transform 1 0 9108 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1870_
timestamp 1644511149
transform 1 0 1748 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1871_
timestamp 1644511149
transform 1 0 1840 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1872_
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1873_
timestamp 1644511149
transform 1 0 30820 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1874_
timestamp 1644511149
transform 1 0 16836 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1875_
timestamp 1644511149
transform 1 0 2116 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1876_
timestamp 1644511149
transform 1 0 31280 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1877_
timestamp 1644511149
transform 1 0 5152 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1878_
timestamp 1644511149
transform 1 0 46276 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1879_
timestamp 1644511149
transform 1 0 23368 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1880_
timestamp 1644511149
transform 1 0 12420 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1881_
timestamp 1644511149
transform 1 0 29716 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1882_
timestamp 1644511149
transform 1 0 20240 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1883_
timestamp 1644511149
transform 1 0 42412 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1884_
timestamp 1644511149
transform 1 0 46276 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1885_
timestamp 1644511149
transform 1 0 4508 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1886_
timestamp 1644511149
transform 1 0 41400 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1887_
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1888_
timestamp 1644511149
transform 1 0 1380 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1889_
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1890_
timestamp 1644511149
transform 1 0 20240 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1891_
timestamp 1644511149
transform 1 0 15088 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1892_
timestamp 1644511149
transform 1 0 29716 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1893_
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1894_
timestamp 1644511149
transform 1 0 46276 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1895_
timestamp 1644511149
transform 1 0 29716 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1896_
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1897_
timestamp 1644511149
transform 1 0 22448 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1898_
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1899_
timestamp 1644511149
transform 1 0 46276 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1900_
timestamp 1644511149
transform 1 0 1932 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1901_
timestamp 1644511149
transform 1 0 46276 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1902_
timestamp 1644511149
transform 1 0 46000 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1903_
timestamp 1644511149
transform 1 0 46276 0 1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1904_
timestamp 1644511149
transform 1 0 1380 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1905_
timestamp 1644511149
transform 1 0 11408 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1906_
timestamp 1644511149
transform 1 0 35604 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1907_
timestamp 1644511149
transform 1 0 35144 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1908_
timestamp 1644511149
transform 1 0 35512 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1909_
timestamp 1644511149
transform 1 0 35512 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1910_
timestamp 1644511149
transform 1 0 35512 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1911_
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1912_
timestamp 1644511149
transform 1 0 7360 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1913_
timestamp 1644511149
transform 1 0 35420 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1914_
timestamp 1644511149
transform 1 0 12420 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1915_
timestamp 1644511149
transform 1 0 46276 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1916_
timestamp 1644511149
transform 1 0 45172 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1917_
timestamp 1644511149
transform 1 0 39192 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1918_
timestamp 1644511149
transform 1 0 9844 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1919_
timestamp 1644511149
transform 1 0 6532 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1920_
timestamp 1644511149
transform 1 0 46276 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1921_
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1922_
timestamp 1644511149
transform 1 0 32292 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1923_
timestamp 1644511149
transform 1 0 34316 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1924_
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1925_
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1926_
timestamp 1644511149
transform 1 0 34500 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1927_
timestamp 1644511149
transform 1 0 34500 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1928_
timestamp 1644511149
transform 1 0 32936 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1929_
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1930_
timestamp 1644511149
transform 1 0 24932 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1931_
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1932_
timestamp 1644511149
transform 1 0 33396 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1933_
timestamp 1644511149
transform 1 0 10856 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1934_
timestamp 1644511149
transform 1 0 6348 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1935_
timestamp 1644511149
transform 1 0 33488 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1936_
timestamp 1644511149
transform 1 0 14444 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1937_
timestamp 1644511149
transform 1 0 1748 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1938_
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1939_
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1940_
timestamp 1644511149
transform 1 0 46276 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1941_
timestamp 1644511149
transform 1 0 44068 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1942_
timestamp 1644511149
transform 1 0 2116 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1943_
timestamp 1644511149
transform 1 0 27968 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1944_
timestamp 1644511149
transform 1 0 46276 0 1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1945_
timestamp 1644511149
transform 1 0 41860 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1946_
timestamp 1644511149
transform 1 0 46276 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1947_
timestamp 1644511149
transform 1 0 3956 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1948_
timestamp 1644511149
transform 1 0 13156 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1949_
timestamp 1644511149
transform 1 0 26680 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1950_
timestamp 1644511149
transform 1 0 42872 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1951_
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1952_
timestamp 1644511149
transform 1 0 42596 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1953_
timestamp 1644511149
transform 1 0 1656 0 -1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1954_
timestamp 1644511149
transform 1 0 46276 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1955_
timestamp 1644511149
transform 1 0 1380 0 1 44608
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1956_
timestamp 1644511149
transform 1 0 46276 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1957_
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1958_
timestamp 1644511149
transform 1 0 46276 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1959_
timestamp 1644511149
transform 1 0 46276 0 1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1960_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1961_
timestamp 1644511149
transform 1 0 46276 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1962_
timestamp 1644511149
transform 1 0 44712 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1963_
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1964_
timestamp 1644511149
transform 1 0 45172 0 1 2176
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1965_
timestamp 1644511149
transform 1 0 8924 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1966_
timestamp 1644511149
transform 1 0 46276 0 1 42432
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1967_
timestamp 1644511149
transform 1 0 46276 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1968_
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1969_
timestamp 1644511149
transform 1 0 1380 0 1 41344
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1970_
timestamp 1644511149
transform 1 0 36064 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1971_
timestamp 1644511149
transform 1 0 45172 0 -1 45696
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1972_
timestamp 1644511149
transform 1 0 1380 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1973_
timestamp 1644511149
transform 1 0 44988 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1974_
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1975_
timestamp 1644511149
transform 1 0 45080 0 -1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1976_
timestamp 1644511149
transform 1 0 24380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1977_
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1978_
timestamp 1644511149
transform 1 0 46276 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1979_
timestamp 1644511149
transform 1 0 1380 0 1 47872
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1980_
timestamp 1644511149
transform 1 0 11684 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1981_
timestamp 1644511149
transform 1 0 45172 0 -1 46784
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1982_
timestamp 1644511149
transform 1 0 1380 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1983_
timestamp 1644511149
transform 1 0 32108 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1984_
timestamp 1644511149
transform 1 0 21804 0 1 48960
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1985_
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1986_
timestamp 1644511149
transform 1 0 1748 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1987_
timestamp 1644511149
transform 1 0 38548 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__ebufn_8  _1988_
timestamp 1644511149
transform 1 0 2024 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_wb_clk_i
timestamp 1644511149
transform 1 0 21620 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 22724 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_1_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 20976 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 26496 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 18308 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_2_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 17296 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 27508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 27876 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 16928 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 17112 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 27600 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_3_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_0_0_wb_clk_i
timestamp 1644511149
transform 1 0 20056 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_1_0_wb_clk_i
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_2_0_wb_clk_i
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_3_0_wb_clk_i
timestamp 1644511149
transform 1 0 18584 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_4_0_wb_clk_i
timestamp 1644511149
transform 1 0 25944 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_5_0_wb_clk_i
timestamp 1644511149
transform 1 0 28888 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_6_0_wb_clk_i
timestamp 1644511149
transform 1 0 27692 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_7_0_wb_clk_i
timestamp 1644511149
transform 1 0 29900 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_8_0_wb_clk_i
timestamp 1644511149
transform 1 0 14904 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_9_0_wb_clk_i
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_10_0_wb_clk_i
timestamp 1644511149
transform 1 0 15364 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_11_0_wb_clk_i
timestamp 1644511149
transform 1 0 20424 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_12_0_wb_clk_i
timestamp 1644511149
transform 1 0 26956 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_13_0_wb_clk_i
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_14_0_wb_clk_i
timestamp 1644511149
transform 1 0 24656 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  clkbuf_4_15_0_wb_clk_i
timestamp 1644511149
transform 1 0 27600 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkdlybuf4s50_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20608 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__buf_6  input1
timestamp 1644511149
transform 1 0 47380 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input2
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform 1 0 14444 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1644511149
transform 1 0 22632 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input6
timestamp 1644511149
transform 1 0 47656 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input7
timestamp 1644511149
transform 1 0 47840 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1644511149
transform 1 0 21068 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input9
timestamp 1644511149
transform 1 0 12696 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1644511149
transform 1 0 18952 0 -1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input11
timestamp 1644511149
transform 1 0 27048 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input12
timestamp 1644511149
transform 1 0 32936 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input13
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input14
timestamp 1644511149
transform 1 0 10212 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input15
timestamp 1644511149
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input16
timestamp 1644511149
transform 1 0 16652 0 1 48960
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input17
timestamp 1644511149
transform 1 0 47656 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1644511149
transform 1 0 47840 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input20
timestamp 1644511149
transform 1 0 47840 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1644511149
transform 1 0 24380 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input22
timestamp 1644511149
transform 1 0 1380 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input23
timestamp 1644511149
transform 1 0 2668 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 47840 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input25
timestamp 1644511149
transform 1 0 1380 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input26
timestamp 1644511149
transform 1 0 47656 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1644511149
transform 1 0 15180 0 1 48960
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1644511149
transform 1 0 47288 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input29
timestamp 1644511149
transform 1 0 47840 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input30
timestamp 1644511149
transform 1 0 3772 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input31
timestamp 1644511149
transform 1 0 5060 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform 1 0 20056 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input33
timestamp 1644511149
transform 1 0 1748 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input34
timestamp 1644511149
transform 1 0 40664 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 27324 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input36
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input37
timestamp 1644511149
transform 1 0 38088 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input38
timestamp 1644511149
transform 1 0 20056 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input40
timestamp 1644511149
transform 1 0 5520 0 -1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input41
timestamp 1644511149
transform 1 0 47840 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform 1 0 1748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input43
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input44
timestamp 1644511149
transform 1 0 1748 0 -1 44608
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input45
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input46
timestamp 1644511149
transform 1 0 43240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 44988 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input48
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1644511149
transform 1 0 25852 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input51
timestamp 1644511149
transform 1 0 47840 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input52
timestamp 1644511149
transform 1 0 19320 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 24564 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input55
timestamp 1644511149
transform 1 0 28704 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1644511149
transform 1 0 47932 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input57
timestamp 1644511149
transform 1 0 47288 0 1 40256
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input58
timestamp 1644511149
transform 1 0 17480 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input59
timestamp 1644511149
transform 1 0 47840 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input60
timestamp 1644511149
transform 1 0 46828 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input61
timestamp 1644511149
transform 1 0 34868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input62
timestamp 1644511149
transform 1 0 47656 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 33856 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input64
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input65
timestamp 1644511149
transform 1 0 1380 0 1 45696
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input66
timestamp 1644511149
transform 1 0 44160 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input67
timestamp 1644511149
transform 1 0 47840 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input68
timestamp 1644511149
transform 1 0 25852 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input69
timestamp 1644511149
transform 1 0 47840 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input70
timestamp 1644511149
transform 1 0 1748 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input71
timestamp 1644511149
transform 1 0 4140 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input72
timestamp 1644511149
transform 1 0 2024 0 -1 46784
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input73
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input74
timestamp 1644511149
transform 1 0 9936 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input75
timestamp 1644511149
transform 1 0 47840 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input76
timestamp 1644511149
transform 1 0 1380 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  input77
timestamp 1644511149
transform 1 0 41400 0 1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input78
timestamp 1644511149
transform 1 0 47656 0 -1 48960
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input79
timestamp 1644511149
transform 1 0 11868 0 1 48960
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input80
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input81
timestamp 1644511149
transform 1 0 47840 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input82
timestamp 1644511149
transform 1 0 47656 0 -1 47872
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1644511149
transform 1 0 1748 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input84
timestamp 1644511149
transform 1 0 47840 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input85
timestamp 1644511149
transform 1 0 1380 0 -1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input86
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input87
timestamp 1644511149
transform 1 0 47840 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1644511149
transform 1 0 22632 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1644511149
transform 1 0 47288 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input91
timestamp 1644511149
transform 1 0 43884 0 1 47872
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input92
timestamp 1644511149
transform 1 0 47840 0 1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input93
timestamp 1644511149
transform 1 0 47840 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input94
timestamp 1644511149
transform 1 0 1748 0 1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input95
timestamp 1644511149
transform 1 0 47840 0 1 25024
box -38 -48 406 592
<< labels >>
rlabel metal3 s 49200 31968 50000 32088 6 active
port 0 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 1368 800 1488 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 38768 800 38888 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 25134 51200 25190 52000 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 49200 15648 50000 15768 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 21270 51200 21326 52000 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 49200 2048 50000 2168 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 io_in[16]
port 8 nsew signal input
rlabel metal3 s 0 14968 800 15088 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 io_in[18]
port 10 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 io_in[1]
port 12 nsew signal input
rlabel metal3 s 49200 18368 50000 18488 6 io_in[20]
port 13 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 49200 21088 50000 21208 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 49200 32648 50000 32768 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 49200 23128 50000 23248 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 2594 51200 2650 52000 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 28998 0 29054 800 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 46386 51200 46442 52000 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 16762 0 16818 800 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 9034 51200 9090 52000 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 31574 51200 31630 52000 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 49200 47608 50000 47728 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 49200 20408 50000 20528 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 35438 51200 35494 52000 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 49200 2728 50000 2848 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 3882 51200 3938 52000 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 0 42848 800 42968 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 io_oeb[0]
port 39 nsew signal tristate
rlabel metal3 s 49200 24488 50000 24608 6 io_oeb[10]
port 40 nsew signal tristate
rlabel metal2 s 45098 0 45154 800 6 io_oeb[11]
port 41 nsew signal tristate
rlabel metal2 s 5814 0 5870 800 6 io_oeb[12]
port 42 nsew signal tristate
rlabel metal2 s 48318 0 48374 800 6 io_oeb[13]
port 43 nsew signal tristate
rlabel metal2 s 7746 51200 7802 52000 6 io_oeb[14]
port 44 nsew signal tristate
rlabel metal3 s 49200 43528 50000 43648 6 io_oeb[15]
port 45 nsew signal tristate
rlabel metal3 s 49200 4768 50000 4888 6 io_oeb[16]
port 46 nsew signal tristate
rlabel metal3 s 0 6808 800 6928 6 io_oeb[17]
port 47 nsew signal tristate
rlabel metal3 s 0 41488 800 41608 6 io_oeb[18]
port 48 nsew signal tristate
rlabel metal2 s 36726 0 36782 800 6 io_oeb[19]
port 49 nsew signal tristate
rlabel metal2 s 43166 51200 43222 52000 6 io_oeb[1]
port 50 nsew signal tristate
rlabel metal3 s 49200 46928 50000 47048 6 io_oeb[20]
port 51 nsew signal tristate
rlabel metal3 s 0 9528 800 9648 6 io_oeb[21]
port 52 nsew signal tristate
rlabel metal2 s 45098 51200 45154 52000 6 io_oeb[22]
port 53 nsew signal tristate
rlabel metal3 s 0 26528 800 26648 6 io_oeb[23]
port 54 nsew signal tristate
rlabel metal3 s 49200 51688 50000 51808 6 io_oeb[24]
port 55 nsew signal tristate
rlabel metal2 s 24490 51200 24546 52000 6 io_oeb[25]
port 56 nsew signal tristate
rlabel metal3 s 0 23128 800 23248 6 io_oeb[26]
port 57 nsew signal tristate
rlabel metal3 s 49200 28568 50000 28688 6 io_oeb[27]
port 58 nsew signal tristate
rlabel metal2 s 1306 51200 1362 52000 6 io_oeb[28]
port 59 nsew signal tristate
rlabel metal2 s 12254 0 12310 800 6 io_oeb[29]
port 60 nsew signal tristate
rlabel metal3 s 0 51688 800 51808 6 io_oeb[2]
port 61 nsew signal tristate
rlabel metal2 s 49606 51200 49662 52000 6 io_oeb[30]
port 62 nsew signal tristate
rlabel metal3 s 0 3408 800 3528 6 io_oeb[31]
port 63 nsew signal tristate
rlabel metal2 s 33506 0 33562 800 6 io_oeb[32]
port 64 nsew signal tristate
rlabel metal2 s 22558 51200 22614 52000 6 io_oeb[33]
port 65 nsew signal tristate
rlabel metal3 s 0 17688 800 17808 6 io_oeb[34]
port 66 nsew signal tristate
rlabel metal3 s 0 13608 800 13728 6 io_oeb[35]
port 67 nsew signal tristate
rlabel metal2 s 39946 0 40002 800 6 io_oeb[36]
port 68 nsew signal tristate
rlabel metal3 s 0 39448 800 39568 6 io_oeb[37]
port 69 nsew signal tristate
rlabel metal3 s 49200 45568 50000 45688 6 io_oeb[3]
port 70 nsew signal tristate
rlabel metal3 s 0 44888 800 45008 6 io_oeb[4]
port 71 nsew signal tristate
rlabel metal3 s 49200 36728 50000 36848 6 io_oeb[5]
port 72 nsew signal tristate
rlabel metal2 s 21270 0 21326 800 6 io_oeb[6]
port 73 nsew signal tristate
rlabel metal3 s 49200 17008 50000 17128 6 io_oeb[7]
port 74 nsew signal tristate
rlabel metal3 s 49200 49648 50000 49768 6 io_oeb[8]
port 75 nsew signal tristate
rlabel metal3 s 49200 16328 50000 16448 6 io_oeb[9]
port 76 nsew signal tristate
rlabel metal2 s 36082 51200 36138 52000 6 io_out[0]
port 77 nsew signal tristate
rlabel metal3 s 49200 44208 50000 44328 6 io_out[10]
port 78 nsew signal tristate
rlabel metal3 s 49200 9528 50000 9648 6 io_out[11]
port 79 nsew signal tristate
rlabel metal2 s 48962 0 49018 800 6 io_out[12]
port 80 nsew signal tristate
rlabel metal2 s 47030 0 47086 800 6 io_out[13]
port 81 nsew signal tristate
rlabel metal3 s 49200 12248 50000 12368 6 io_out[14]
port 82 nsew signal tristate
rlabel metal2 s 37370 0 37426 800 6 io_out[15]
port 83 nsew signal tristate
rlabel metal2 s 37370 51200 37426 52000 6 io_out[16]
port 84 nsew signal tristate
rlabel metal2 s 38658 51200 38714 52000 6 io_out[17]
port 85 nsew signal tristate
rlabel metal2 s 15474 51200 15530 52000 6 io_out[18]
port 86 nsew signal tristate
rlabel metal3 s 49200 3408 50000 3528 6 io_out[19]
port 87 nsew signal tristate
rlabel metal2 s 12898 0 12954 800 6 io_out[1]
port 88 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 io_out[20]
port 89 nsew signal tristate
rlabel metal3 s 0 48288 800 48408 6 io_out[21]
port 90 nsew signal tristate
rlabel metal2 s 34794 51200 34850 52000 6 io_out[22]
port 91 nsew signal tristate
rlabel metal2 s 14830 51200 14886 52000 6 io_out[23]
port 92 nsew signal tristate
rlabel metal3 s 0 46248 800 46368 6 io_out[24]
port 93 nsew signal tristate
rlabel metal3 s 0 34008 800 34128 6 io_out[25]
port 94 nsew signal tristate
rlabel metal3 s 0 27208 800 27328 6 io_out[26]
port 95 nsew signal tristate
rlabel metal3 s 49200 7488 50000 7608 6 io_out[27]
port 96 nsew signal tristate
rlabel metal2 s 44454 0 44510 800 6 io_out[28]
port 97 nsew signal tristate
rlabel metal3 s 0 5448 800 5568 6 io_out[29]
port 98 nsew signal tristate
rlabel metal3 s 49200 35368 50000 35488 6 io_out[2]
port 99 nsew signal tristate
rlabel metal2 s 28354 51200 28410 52000 6 io_out[30]
port 100 nsew signal tristate
rlabel metal3 s 49200 46248 50000 46368 6 io_out[31]
port 101 nsew signal tristate
rlabel metal2 s 42522 0 42578 800 6 io_out[32]
port 102 nsew signal tristate
rlabel metal3 s 49200 10888 50000 11008 6 io_out[33]
port 103 nsew signal tristate
rlabel metal3 s 0 51008 800 51128 6 io_out[34]
port 104 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 io_out[35]
port 105 nsew signal tristate
rlabel metal2 s 27066 51200 27122 52000 6 io_out[36]
port 106 nsew signal tristate
rlabel metal2 s 48318 51200 48374 52000 6 io_out[37]
port 107 nsew signal tristate
rlabel metal2 s 45742 51200 45798 52000 6 io_out[3]
port 108 nsew signal tristate
rlabel metal2 s 39946 51200 40002 52000 6 io_out[4]
port 109 nsew signal tristate
rlabel metal2 s 10322 51200 10378 52000 6 io_out[5]
port 110 nsew signal tristate
rlabel metal2 s 7102 51200 7158 52000 6 io_out[6]
port 111 nsew signal tristate
rlabel metal3 s 49200 34008 50000 34128 6 io_out[7]
port 112 nsew signal tristate
rlabel metal2 s 2594 0 2650 800 6 io_out[8]
port 113 nsew signal tristate
rlabel metal2 s 8390 51200 8446 52000 6 io_out[9]
port 114 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 rambus_wb_ack_i
port 115 nsew signal input
rlabel metal3 s 49200 40128 50000 40248 6 rambus_wb_adr_o[0]
port 116 nsew signal tristate
rlabel metal3 s 0 46928 800 47048 6 rambus_wb_adr_o[1]
port 117 nsew signal tristate
rlabel metal2 s 10966 51200 11022 52000 6 rambus_wb_adr_o[2]
port 118 nsew signal tristate
rlabel metal3 s 49200 6128 50000 6248 6 rambus_wb_adr_o[3]
port 119 nsew signal tristate
rlabel metal3 s 49200 51008 50000 51128 6 rambus_wb_adr_o[4]
port 120 nsew signal tristate
rlabel metal3 s 49200 17688 50000 17808 6 rambus_wb_adr_o[5]
port 121 nsew signal tristate
rlabel metal3 s 49200 6808 50000 6928 6 rambus_wb_adr_o[6]
port 122 nsew signal tristate
rlabel metal3 s 49200 29248 50000 29368 6 rambus_wb_adr_o[7]
port 123 nsew signal tristate
rlabel metal2 s 9034 0 9090 800 6 rambus_wb_adr_o[8]
port 124 nsew signal tristate
rlabel metal3 s 0 2048 800 2168 6 rambus_wb_adr_o[9]
port 125 nsew signal tristate
rlabel metal3 s 0 18368 800 18488 6 rambus_wb_clk_o
port 126 nsew signal tristate
rlabel metal2 s 5170 51200 5226 52000 6 rambus_wb_cyc_o
port 127 nsew signal tristate
rlabel metal2 s 13542 51200 13598 52000 6 rambus_wb_dat_i[0]
port 128 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 rambus_wb_dat_i[10]
port 129 nsew signal input
rlabel metal3 s 0 22448 800 22568 6 rambus_wb_dat_i[11]
port 130 nsew signal input
rlabel metal3 s 49200 688 50000 808 6 rambus_wb_dat_i[12]
port 131 nsew signal input
rlabel metal3 s 49200 13608 50000 13728 6 rambus_wb_dat_i[13]
port 132 nsew signal input
rlabel metal2 s 21914 51200 21970 52000 6 rambus_wb_dat_i[14]
port 133 nsew signal input
rlabel metal2 s 12898 51200 12954 52000 6 rambus_wb_dat_i[15]
port 134 nsew signal input
rlabel metal2 s 18050 51200 18106 52000 6 rambus_wb_dat_i[16]
port 135 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 rambus_wb_dat_i[17]
port 136 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 rambus_wb_dat_i[18]
port 137 nsew signal input
rlabel metal3 s 0 34688 800 34808 6 rambus_wb_dat_i[19]
port 138 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 rambus_wb_dat_i[1]
port 139 nsew signal input
rlabel metal3 s 0 7488 800 7608 6 rambus_wb_dat_i[20]
port 140 nsew signal input
rlabel metal2 s 16118 51200 16174 52000 6 rambus_wb_dat_i[21]
port 141 nsew signal input
rlabel metal3 s 49200 8168 50000 8288 6 rambus_wb_dat_i[22]
port 142 nsew signal input
rlabel metal3 s 49200 31288 50000 31408 6 rambus_wb_dat_i[23]
port 143 nsew signal input
rlabel metal3 s 49200 33328 50000 33448 6 rambus_wb_dat_i[24]
port 144 nsew signal input
rlabel metal3 s 49200 38768 50000 38888 6 rambus_wb_dat_i[25]
port 145 nsew signal input
rlabel metal2 s 23846 51200 23902 52000 6 rambus_wb_dat_i[26]
port 146 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 rambus_wb_dat_i[27]
port 147 nsew signal input
rlabel metal2 s 18 51200 74 52000 6 rambus_wb_dat_i[28]
port 148 nsew signal input
rlabel metal3 s 49200 42168 50000 42288 6 rambus_wb_dat_i[29]
port 149 nsew signal input
rlabel metal3 s 0 40128 800 40248 6 rambus_wb_dat_i[2]
port 150 nsew signal input
rlabel metal3 s 49200 10208 50000 10328 6 rambus_wb_dat_i[30]
port 151 nsew signal input
rlabel metal2 s 14186 51200 14242 52000 6 rambus_wb_dat_i[31]
port 152 nsew signal input
rlabel metal3 s 49200 29928 50000 30048 6 rambus_wb_dat_i[3]
port 153 nsew signal input
rlabel metal3 s 49200 23808 50000 23928 6 rambus_wb_dat_i[4]
port 154 nsew signal input
rlabel metal3 s 0 47608 800 47728 6 rambus_wb_dat_i[5]
port 155 nsew signal input
rlabel metal2 s 4526 51200 4582 52000 6 rambus_wb_dat_i[6]
port 156 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 rambus_wb_dat_i[7]
port 157 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 rambus_wb_dat_i[8]
port 158 nsew signal input
rlabel metal2 s 40590 51200 40646 52000 6 rambus_wb_dat_i[9]
port 159 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 rambus_wb_dat_o[0]
port 160 nsew signal tristate
rlabel metal2 s 30286 0 30342 800 6 rambus_wb_dat_o[10]
port 161 nsew signal tristate
rlabel metal2 s 20626 0 20682 800 6 rambus_wb_dat_o[11]
port 162 nsew signal tristate
rlabel metal2 s 41878 0 41934 800 6 rambus_wb_dat_o[12]
port 163 nsew signal tristate
rlabel metal3 s 49200 34688 50000 34808 6 rambus_wb_dat_o[13]
port 164 nsew signal tristate
rlabel metal3 s 0 50328 800 50448 6 rambus_wb_dat_o[14]
port 165 nsew signal tristate
rlabel metal2 s 42522 51200 42578 52000 6 rambus_wb_dat_o[15]
port 166 nsew signal tristate
rlabel metal2 s 1306 0 1362 800 6 rambus_wb_dat_o[16]
port 167 nsew signal tristate
rlabel metal3 s 0 29928 800 30048 6 rambus_wb_dat_o[17]
port 168 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 rambus_wb_dat_o[18]
port 169 nsew signal tristate
rlabel metal2 s 20626 51200 20682 52000 6 rambus_wb_dat_o[19]
port 170 nsew signal tristate
rlabel metal3 s 0 10208 800 10328 6 rambus_wb_dat_o[1]
port 171 nsew signal tristate
rlabel metal2 s 15474 0 15530 800 6 rambus_wb_dat_o[20]
port 172 nsew signal tristate
rlabel metal2 s 30930 0 30986 800 6 rambus_wb_dat_o[21]
port 173 nsew signal tristate
rlabel metal3 s 0 31968 800 32088 6 rambus_wb_dat_o[22]
port 174 nsew signal tristate
rlabel metal3 s 49200 19728 50000 19848 6 rambus_wb_dat_o[23]
port 175 nsew signal tristate
rlabel metal2 s 30930 51200 30986 52000 6 rambus_wb_dat_o[24]
port 176 nsew signal tristate
rlabel metal3 s 0 16328 800 16448 6 rambus_wb_dat_o[25]
port 177 nsew signal tristate
rlabel metal2 s 23202 51200 23258 52000 6 rambus_wb_dat_o[26]
port 178 nsew signal tristate
rlabel metal3 s 0 28568 800 28688 6 rambus_wb_dat_o[27]
port 179 nsew signal tristate
rlabel metal3 s 49200 50328 50000 50448 6 rambus_wb_dat_o[28]
port 180 nsew signal tristate
rlabel metal3 s 0 48968 800 49088 6 rambus_wb_dat_o[29]
port 181 nsew signal tristate
rlabel metal2 s 31574 0 31630 800 6 rambus_wb_dat_o[2]
port 182 nsew signal tristate
rlabel metal3 s 49200 41488 50000 41608 6 rambus_wb_dat_o[30]
port 183 nsew signal tristate
rlabel metal2 s 46386 0 46442 800 6 rambus_wb_dat_o[31]
port 184 nsew signal tristate
rlabel metal2 s 17406 51200 17462 52000 6 rambus_wb_dat_o[3]
port 185 nsew signal tristate
rlabel metal3 s 0 32648 800 32768 6 rambus_wb_dat_o[4]
port 186 nsew signal tristate
rlabel metal2 s 32218 51200 32274 52000 6 rambus_wb_dat_o[5]
port 187 nsew signal tristate
rlabel metal2 s 5170 0 5226 800 6 rambus_wb_dat_o[6]
port 188 nsew signal tristate
rlabel metal3 s 49200 14288 50000 14408 6 rambus_wb_dat_o[7]
port 189 nsew signal tristate
rlabel metal2 s 23846 0 23902 800 6 rambus_wb_dat_o[8]
port 190 nsew signal tristate
rlabel metal2 s 12254 51200 12310 52000 6 rambus_wb_dat_o[9]
port 191 nsew signal tristate
rlabel metal3 s 0 8848 800 8968 6 rambus_wb_rst_o
port 192 nsew signal tristate
rlabel metal2 s 41234 0 41290 800 6 rambus_wb_sel_o[0]
port 193 nsew signal tristate
rlabel metal2 s 32862 51200 32918 52000 6 rambus_wb_sel_o[1]
port 194 nsew signal tristate
rlabel metal2 s 9678 51200 9734 52000 6 rambus_wb_sel_o[2]
port 195 nsew signal tristate
rlabel metal3 s 0 33328 800 33448 6 rambus_wb_sel_o[3]
port 196 nsew signal tristate
rlabel metal2 s 29642 51200 29698 52000 6 rambus_wb_stb_o
port 197 nsew signal tristate
rlabel metal3 s 0 4768 800 4888 6 rambus_wb_we_o
port 198 nsew signal tristate
rlabel metal4 s 4208 2128 4528 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 34928 2128 35248 49552 6 vccd1
port 199 nsew power input
rlabel metal4 s 19568 2128 19888 49552 6 vssd1
port 200 nsew ground input
rlabel metal3 s 49200 1368 50000 1488 6 wb_clk_i
port 201 nsew signal input
rlabel metal2 s 26422 51200 26478 52000 6 wb_rst_i
port 202 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 wbs_ack_o
port 203 nsew signal tristate
rlabel metal3 s 0 31288 800 31408 6 wbs_adr_i[0]
port 204 nsew signal input
rlabel metal2 s 38014 51200 38070 52000 6 wbs_adr_i[10]
port 205 nsew signal input
rlabel metal2 s 19982 51200 20038 52000 6 wbs_adr_i[11]
port 206 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 wbs_adr_i[12]
port 207 nsew signal input
rlabel metal2 s 6458 51200 6514 52000 6 wbs_adr_i[13]
port 208 nsew signal input
rlabel metal3 s 49200 27888 50000 28008 6 wbs_adr_i[14]
port 209 nsew signal input
rlabel metal3 s 0 688 800 808 6 wbs_adr_i[15]
port 210 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_adr_i[16]
port 211 nsew signal input
rlabel metal3 s 0 44208 800 44328 6 wbs_adr_i[17]
port 212 nsew signal input
rlabel metal3 s 0 17008 800 17128 6 wbs_adr_i[18]
port 213 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 wbs_adr_i[19]
port 214 nsew signal input
rlabel metal2 s 44454 51200 44510 52000 6 wbs_adr_i[1]
port 215 nsew signal input
rlabel metal3 s 0 23808 800 23928 6 wbs_adr_i[20]
port 216 nsew signal input
rlabel metal2 s 25134 0 25190 800 6 wbs_adr_i[21]
port 217 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 wbs_adr_i[22]
port 218 nsew signal input
rlabel metal3 s 49200 5448 50000 5568 6 wbs_adr_i[23]
port 219 nsew signal input
rlabel metal2 s 19338 51200 19394 52000 6 wbs_adr_i[24]
port 220 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 wbs_adr_i[25]
port 221 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_adr_i[26]
port 222 nsew signal input
rlabel metal2 s 28998 51200 29054 52000 6 wbs_adr_i[27]
port 223 nsew signal input
rlabel metal3 s 49200 22448 50000 22568 6 wbs_adr_i[28]
port 224 nsew signal input
rlabel metal3 s 49200 40808 50000 40928 6 wbs_adr_i[29]
port 225 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[2]
port 226 nsew signal input
rlabel metal2 s 48962 51200 49018 52000 6 wbs_adr_i[30]
port 227 nsew signal input
rlabel metal3 s 49200 14968 50000 15088 6 wbs_adr_i[31]
port 228 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 wbs_adr_i[3]
port 229 nsew signal input
rlabel metal2 s 47674 51200 47730 52000 6 wbs_adr_i[4]
port 230 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 wbs_adr_i[5]
port 231 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_adr_i[6]
port 232 nsew signal input
rlabel metal3 s 0 45568 800 45688 6 wbs_adr_i[7]
port 233 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 wbs_adr_i[8]
port 234 nsew signal input
rlabel metal3 s 49200 8848 50000 8968 6 wbs_adr_i[9]
port 235 nsew signal input
rlabel metal2 s 25778 51200 25834 52000 6 wbs_cyc_i
port 236 nsew signal input
rlabel metal3 s 49200 38088 50000 38208 6 wbs_dat_i[0]
port 237 nsew signal input
rlabel metal2 s 662 51200 718 52000 6 wbs_dat_i[10]
port 238 nsew signal input
rlabel metal2 s 3238 51200 3294 52000 6 wbs_dat_i[11]
port 239 nsew signal input
rlabel metal2 s 1950 51200 2006 52000 6 wbs_dat_i[12]
port 240 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[13]
port 241 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[14]
port 242 nsew signal input
rlabel metal3 s 49200 21768 50000 21888 6 wbs_dat_i[15]
port 243 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 wbs_dat_i[16]
port 244 nsew signal input
rlabel metal2 s 41878 51200 41934 52000 6 wbs_dat_i[17]
port 245 nsew signal input
rlabel metal3 s 49200 48968 50000 49088 6 wbs_dat_i[18]
port 246 nsew signal input
rlabel metal2 s 11610 51200 11666 52000 6 wbs_dat_i[19]
port 247 nsew signal input
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_i[1]
port 248 nsew signal input
rlabel metal3 s 49200 25848 50000 25968 6 wbs_dat_i[20]
port 249 nsew signal input
rlabel metal3 s 49200 48288 50000 48408 6 wbs_dat_i[21]
port 250 nsew signal input
rlabel metal3 s 0 40808 800 40928 6 wbs_dat_i[22]
port 251 nsew signal input
rlabel metal3 s 49200 36048 50000 36168 6 wbs_dat_i[23]
port 252 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 wbs_dat_i[24]
port 253 nsew signal input
rlabel metal3 s 0 15648 800 15768 6 wbs_dat_i[25]
port 254 nsew signal input
rlabel metal2 s 47030 51200 47086 52000 6 wbs_dat_i[26]
port 255 nsew signal input
rlabel metal2 s 18694 51200 18750 52000 6 wbs_dat_i[27]
port 256 nsew signal input
rlabel metal2 s 14830 0 14886 800 6 wbs_dat_i[28]
port 257 nsew signal input
rlabel metal3 s 49200 27208 50000 27328 6 wbs_dat_i[29]
port 258 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 wbs_dat_i[2]
port 259 nsew signal input
rlabel metal3 s 49200 11568 50000 11688 6 wbs_dat_i[30]
port 260 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 wbs_dat_i[31]
port 261 nsew signal input
rlabel metal2 s 49606 0 49662 800 6 wbs_dat_i[3]
port 262 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[4]
port 263 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 wbs_dat_i[5]
port 264 nsew signal input
rlabel metal3 s 49200 19048 50000 19168 6 wbs_dat_i[6]
port 265 nsew signal input
rlabel metal2 s 43810 51200 43866 52000 6 wbs_dat_i[7]
port 266 nsew signal input
rlabel metal3 s 49200 42848 50000 42968 6 wbs_dat_i[8]
port 267 nsew signal input
rlabel metal3 s 49200 8 50000 128 6 wbs_dat_i[9]
port 268 nsew signal input
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[0]
port 269 nsew signal tristate
rlabel metal3 s 49200 26528 50000 26648 6 wbs_dat_o[10]
port 270 nsew signal tristate
rlabel metal2 s 662 0 718 800 6 wbs_dat_o[11]
port 271 nsew signal tristate
rlabel metal3 s 49200 44888 50000 45008 6 wbs_dat_o[12]
port 272 nsew signal tristate
rlabel metal2 s 41234 51200 41290 52000 6 wbs_dat_o[13]
port 273 nsew signal tristate
rlabel metal3 s 49200 4088 50000 4208 6 wbs_dat_o[14]
port 274 nsew signal tristate
rlabel metal2 s 39302 51200 39358 52000 6 wbs_dat_o[15]
port 275 nsew signal tristate
rlabel metal3 s 0 19728 800 19848 6 wbs_dat_o[16]
port 276 nsew signal tristate
rlabel metal3 s 0 21768 800 21888 6 wbs_dat_o[17]
port 277 nsew signal tristate
rlabel metal2 s 32218 0 32274 800 6 wbs_dat_o[18]
port 278 nsew signal tristate
rlabel metal2 s 18 0 74 800 6 wbs_dat_o[19]
port 279 nsew signal tristate
rlabel metal2 s 38014 0 38070 800 6 wbs_dat_o[1]
port 280 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 wbs_dat_o[20]
port 281 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 wbs_dat_o[21]
port 282 nsew signal tristate
rlabel metal3 s 0 12928 800 13048 6 wbs_dat_o[22]
port 283 nsew signal tristate
rlabel metal3 s 0 21088 800 21208 6 wbs_dat_o[23]
port 284 nsew signal tristate
rlabel metal2 s 10322 0 10378 800 6 wbs_dat_o[24]
port 285 nsew signal tristate
rlabel metal2 s 3238 0 3294 800 6 wbs_dat_o[25]
port 286 nsew signal tristate
rlabel metal2 s 27710 51200 27766 52000 6 wbs_dat_o[26]
port 287 nsew signal tristate
rlabel metal2 s 16762 51200 16818 52000 6 wbs_dat_o[27]
port 288 nsew signal tristate
rlabel metal2 s 26422 0 26478 800 6 wbs_dat_o[28]
port 289 nsew signal tristate
rlabel metal2 s 36726 51200 36782 52000 6 wbs_dat_o[29]
port 290 nsew signal tristate
rlabel metal3 s 49200 12928 50000 13048 6 wbs_dat_o[2]
port 291 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 wbs_dat_o[30]
port 292 nsew signal tristate
rlabel metal3 s 49200 39448 50000 39568 6 wbs_dat_o[31]
port 293 nsew signal tristate
rlabel metal2 s 10966 0 11022 800 6 wbs_dat_o[3]
port 294 nsew signal tristate
rlabel metal2 s 18694 0 18750 800 6 wbs_dat_o[4]
port 295 nsew signal tristate
rlabel metal3 s 0 6128 800 6248 6 wbs_dat_o[5]
port 296 nsew signal tristate
rlabel metal3 s 49200 37408 50000 37528 6 wbs_dat_o[6]
port 297 nsew signal tristate
rlabel metal2 s 29642 0 29698 800 6 wbs_dat_o[7]
port 298 nsew signal tristate
rlabel metal2 s 34150 51200 34206 52000 6 wbs_dat_o[8]
port 299 nsew signal tristate
rlabel metal2 s 33506 51200 33562 52000 6 wbs_dat_o[9]
port 300 nsew signal tristate
rlabel metal3 s 0 49648 800 49768 6 wbs_sel_i[0]
port 301 nsew signal input
rlabel metal2 s 5814 51200 5870 52000 6 wbs_sel_i[1]
port 302 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 wbs_sel_i[2]
port 303 nsew signal input
rlabel metal3 s 0 11568 800 11688 6 wbs_sel_i[3]
port 304 nsew signal input
rlabel metal3 s 0 43528 800 43648 6 wbs_stb_i
port 305 nsew signal input
rlabel metal3 s 49200 25168 50000 25288 6 wbs_we_i
port 306 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 50000 52000
<< end >>
